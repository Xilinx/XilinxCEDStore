`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
tIa+y/whfzug+PmRB8SZeZ5chCt3h6t3jKITWLPyiDMx/uTHrOJTPUmHcGuia9oCwh8jq6xOgFco
JKyv+LjDgNXz5ktNhCXca2eA0vylEbcFmqh6Pdo5bphd8L+CYogiUnfF4wNLIHWnpt/0kDyAnzK7
NJv3P0ul7xPXS+Ic+cd5THR5DdBzQjfvu9Dk99HKsaQ/QVdpemmyDrmoTb1KH5DDqx6aDUHQOatX
w71vf1bYGALcd0UD3SMAtNmYaSupWw9y8O6wj7mSC7VzMrk4VBR/C9rGv4xkuygxjHTfj1XR/Uij
BAMLozNLnWrANRFWodFSSnk0n3qVuxKu2xTotw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
okJiP2M+IRsd5WZKqF0Oc8tUEAz7LdKWyebeksLFK8KRBSNGby71R6DD+pTv0OuwTYPsl/0/ADOd
hHVuwJeO9zJFocqw1mwjr3WWzksRCeiJOIplkWcPPYfipYrWaIQOIcdsidKfnmokV4bAUqs5FmSo
TkZImtkxp808vst6BMtDIhAvFHB4zIo2txfih+/G/Vkh5pbs3aJfUTLUG+TEdlvEKLTgy+pVs/Ui
lFU6Rq06BDZ+l4zROHEr3SUJEiFrOd3Y30Qzn66FYUsLp+061Ej/AHe+NiG7+waw3EB7t0SGWEAP
Q4L35V52KOt7ZPfG5rlbnEoRMDf6Wz4ruyYVgQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
TyRBGMva2BLBESRrcH6cdmApxY+ZoiTUtU+ByHbz76sxvvudcmaAt5dvxLsobS9gGUJjaYcF3IBh
g8veVjLayGZTcweVM9BiECKaDyPoTJd2rZScAy9nh8kQiwU6UAIiPV+j3tqr+COvcY+xlJp4doQA
3s4SG3I1dT6bz+s4TeY=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
9Y5bIlwzndHqj1dNiyQRl9EvyN+YvjfaYsNFFCCBIs8W+xnqt38Mm90nQ0iuob3k8bb0/E4SfgIU
l3Sk/0y2ZOF8bF5fLvYKVxzNV5w9z9bq6lnmHbD3B4UHRmFQUVenETD+IDh4OiTmh9wt9HoLQrhU
fcr420COu7Tt0MW9olEJmc0DUQ33T6Nw+uv4ziCG5JOy5X8KLTmV2kCXs5ZM3TcZVEH5FKIB53KS
3s8bsy3+a4XxjVKRfVC4+DZZ8HF58zxL2BZRTa0594vvvtNmoaQVWH0xq6RHauw20uRbzV+KVJAK
Cxm1gsBr1XEAJr5o1axBfz9iJv3JBMPYXbogulktpe7zadcd1WwhJY43vIfHh0mqfyQVFJ4liJww
SNQKApaKZ+zj6YKrfx8bdghZASK2TS747IPvPg6dTJl7nk2+hz8HoCoiN9Y/PJQ3zXbXPp/Y+jK8
xlvnJZDXMLOJYBJAAGLU28GX5aOSaXW9zVh77eVJPgaHER2Lm1b960D1wDATknLks7oIv5vARpCi
7lYgp6gQEDjgzQu1JCKFQMZ4+rUn0c1w927lkEXWgUGtlb3crw/B27HMgXJSrMX1FMr7Fi0mrKRW
Ov/KxcBMxFra10prMhTG5WD1H8UhHxH6/wE5IB28EkFqgdl6iPEK1t/kU13ehjI/NskO5mLLFvbX
NiK2L68fZJY+YajhvSZ9lkwbzW2tktCImN2qh9aGNiJ9cYTvrrrFAV7ONlVx7LxeuJGFo9WO0BSv
CKNzG7L3MsTxGvidiSwKGZrhM3FCZtEZVNWtyzxKE0hpu9NJChyY/gasZs1X0swYFWE77MTmSwbA
02JIFii2o3ycnOnaC7ASuwbAZJgNrAGZ9IR2xnuQ/DKclZ3KYPK7cVu8taWF5CwEXOmH68SSZrNg
Gl/7aoKVaHBvX6bk6uRbWDbGQiz+g/WINm03Psm3HE4+b91cnl+Q3aQ3F+bMz9M+4dNNxjt+4M6+
lIJL65UFJuHNKC0k9Tlu1gdYEdg+m381vpzXiKTVXEvaatKAAeEDPq0nb3yi+Uu7wICIz0jyqrbk
6HGHGWDLWtmYcb1VxfEEDFY1/gA+qCV1kw9cs4qfrbbYiLJMZIzNU7Xwai9UoUjbJzZzwyN8rb57
DwdbjGsI+Hv0Ly4TRXCJAE25+cS3LWFdj8HylR42pK0T66KMXsl1Sklk2YXOqewH3buCGRCJElc4
tmMMDSJPjkwv/igMn/niINDykuW7XxEhfSPLnIgl3L+Xj4rGGWRk8SKk/HE702Rxbv7JgQ/+tZIk
kcvR/06ZwMwR1pnlnMNuXTW5u0W3monQqhIfuA/2uak6rHvPgQFOSqxQ2vJUsoriZRCIbtABWLPH
e+76OqS+sY5QPW/Ok+gnOsuO7DKMeq1rYu+jrvuFYHPXcw4/agz6ESODLW83TXtjWJKuvfFtAqfF
9em1CFDn194TPDyLMd9twHyaST2IPZoAHqTlwTs76HBfsGkhqIzNkvzw8pnwHSj+B4EnjcRHYcFS
whEes5OxG020xV6svBboMcQirAkikbtsctycgKrfjGH3XIU4THQGlIYbgbsOo4u6qTBhCtpTgyaE
Fs5/dLFzvHMxYNvCMJwGwxsZ1k1Zak6nr3KEP/iuCzQ1qm7pdxwfk588pXh5ufrn2Fk8TEAKI9IN
JAheL1uHyTvw3GHTOmeS6vFAEgqdHpul8tRcbW3L848KdDVTUs+zQmHkNd5BaBNGrfDh8eRA8RhP
Upajq1iPgWa3tY2xjPanWqKkH7dUAiZoBKiXT+QhlIP9wE/VgClBvztPYS8YBkBX+6q4PcTbiR79
HtvpTVJkZxRtYxf0EaAV4OpV9CEyUHfa4T5WzS5x7UhLKvYUC1ZxOEc15vshlhtziTCvcOybczuf
F98jkNovfejDumDdvN3hTW0kca7pWJjaCfziMVkohyN2PqlmPgHTGrpii2WAA+7uEKZ1pcq53L8K
cF6JJ4mmdcWg2jcKG7Zmh3sD+ecyQRLVBFeKn2LIb+eAZMPLUTiIlNoJqN1ua8gM469p4C0Qu15h
lPR1QtPEX+4y+TeAaTU/7pq3xCEQwQ8C7n5nmDZimCdDQLUEKOziUe3LMmuGV7Dl17RAn3UYDn3X
Oh/fTscsH09PYQSWhLf5fDUZfa2EC80vmyfRyLiatyTP+vxI8ymTcZxrSIzvD6anwhPfOIy4qxfo
fvVLqMu2AfojMKkWmN0e9C+8yDdXRMWYLuJZ0lyIzK9uUoRGAMRS7/Ws21YptewKbh474JYSaz/T
Djid/I0DrK4Ik74xQRqWo1BqFTka15UiIkEP/lNBObDtQo59dy/4+JDOY/Nh6jnzaOAggqIufUfP
AjUvyBafg2lHh70X9f8bkzq0g/7fa7COoAABlGlEIxm3jvyGc73B2I9BhpyxNOWtYls6J9xtGaNM
IB4qAzFNBkMROR/rNV3SzW34I32iJpbJLT2hRjPz7fjQUS3Zu0iDG5Y/GJSE+GfEmMPZgh6gXBir
PBHDHWwjtlW3qk3sLEKu/KteUsFSWWVnc1riFOhMdNnmFunwORNqgsBgGjiRjugXLG8oyktKsd4A
8kyapU1R0wUJOJwBMn0uuoMSh++Gf9MxhOalZ8bbUSovv+05aUC5lar9D8BUFNW3YxfUISTsK9OJ
+two79tkL1yNLY8+nU+V1lRdK0hyDiW/GsyYtRWi2i9ZSTebjoSRE1cN89ba6eJ6Kr4VOv+iu6ri
5gtfnkM1CFfd7POnyzvJ6Snl38NVia5K4WdFL4RLHpuLjC9nXyl+7hm3EtN/A6TTjXNZd1egx+3n
GpNKrxVq7GG1DjxV1QFBRnj34O0XgcrYuPjo6K+CNhQPQnD6EseiD6sdIy1Vlpp7eLcGnz6WA06I
JSIJd3zcvoN2B9wEOjfEBQU7GHg5tfINXQ+FMCKkDv8reRX8K6o+TuVaod0Xkx3cnGB0LlaljxSP
4UVcyurardAMVLfjxxL/b08Obr4hn1CuZy2FGuLKyZTydzWsNQvtQaKDDeAAGoeyUICI71RW5hrW
THorUYsf6Tg4cI7/4NBkTJC7es+Qs3/fR0RgXAsZQPp3Q1HUHxjyAWKozPbwU2J0/tIzUeRBNSyy
qYbenl5ZdUxIoevffNcWEm7NVB6LIzZPwrWjVND/Ay+eYSQtmN4dbygtfVwYeMUDzYFXofED1U/m
voLSuEwS7T9f03ip2fi6zO5xd8gIcNwE+exXyJHlHn3pQY4k8yjmvr2UBpHh0epVdlEVC3Pnc0Rp
GcyzydOEzCWw0jVFb19PbbpzoNattHc1XsaMRWk4nJjsBfPiKI/nA4ILVM5I0UG/n78S6ziqWbA2
I9m8SncQK3I9LM5VFnbmwtp18zxE9RVwzfP0G7UA7x4mDHVL0uBX6bUZcI/ZQ8rZzcD+cH1ZZy+P
xYCibvVxg6DBWWYiCGD85R+hmxCTWdZqwpY8DfeFkiYzPxdPYgNyuarzhwzxcvnUM2xZAg3ZEycj
waKiN9mErMLi7aTYdJYsrmPTskRLMKSgfhUmSx5IA18BbihWCvUvu/WHODVl+320s/jqr8KiaFe/
K39xUNQWR5akuOEbQrPQS56X90gl2kLJafEdLEYcn5NbRo60sn56QzakDNJ0jYLg5tQ+6CtEj6j/
nbQbmo5Z9Os9FSylrlPEhBdQX5cBBprWry4wiYZDOMlhP/4ARKAo/XZcW4O0y2JfgeHo9vSO0a9Y
niS3BCWx9sFIDPvaM1j8+YWbDTbF8ZAQsyYXptOA+wxIt20PhW4b6umBmERx+wmSpMoMbiA81ggQ
QaI+mjlhpEv8g772yb3sxHJIKFntWK8gMtbm4fX8vUoblaoQoavg4uF44GgNFSWeYNWaVM4oP8RR
LxYvnyRigJu0c3zpsDCLGw6OeF35b4vqLTh2E9DMJFtND1o3pURPt5LzRf5M4CGsGjIJKiydcnjT
q1NQt0Nr2QqaqnPSEK31Z40wUW3op99K9TFYmuNJJsBmDDWbjkQ4ilOKpzeqCEDOwHH2083lALyZ
hlOoYZrYSkFqllW0yufgbs5WWPcGL7lxHrgna+Cz4F9GHrMgAMendmrG1n9kfUTRGSkrcUOSHIg8
IjAiG1xpMqsCjAikwtyfpqC9g7D9TIyirhtuvzgcu+Bg3hiawsKCQTKuz2qSHpuF8gfz/ifxzlwk
N/zWWSGPnZfGvUfCM2Q4lpQthTf/tqeTEEDS1Q8kJEG4g9uVMHXpNLYrpWSHeB6KWJdAgpEdW+/W
3sO8+14s+7+X2O3Zr2p7nhdOG9auVhCWjWBvXb2XqfW8CVExJALqvBJesPibSxWqbpONSPU75+mz
WHdtmOcdlasbezifwisqkhUC/dc5qTIqFPs7X7fB5nrZ/IRUIv40K/z6sfRW4O6WBfU1xK6I7lRq
v4q50FdMt9F/5froMHfFhVo6DGW5TtKCr10vDJGGvRSv5a5n4LJFxlBsds80WNYSDuFmhTc3XYaY
CL7AqJnI/DvbL1Caq0/HolYTDJKBwyzG3RC1uYKVTFjWJ95ftR6M84HQOTDpiAZ6dWpMGEo+Y1bk
9oSLjzN+Lv/TdywK8+YScYzwJWB6KsaifUCQhWhWF40QOJZS1Rtu1cTLcb4tVnxA79fX+b198GFn
JBcbw40TA7sxvOm8CQANriLPkCGB015nc+5RXNy62VtooGNRiAsmw6yE+l9TzTUm3qXFLD2LRfqy
NERq7nTAVXYzd4Ht1O9L1E1vIrFihQvYiysYVXlOwY6nuQWhHnk1dVwHTuJ3/26YbMLHL00s7a0E
s7VCN9PYOSbRm8HPTpIkQcLp8YEpR6BwqPXauAsIYNduYQT998jquYgn/I51QSCZMtLu5hlT9HG0
TjojrTeq+TwSFhH+EZhSQUqWt0tiOxFA0xba1CscjtZy6iRzUo7obGvRg0o2lrsPz/6XZndzbeX+
op1ARXPoPQFbZsDuHGmWjQgN67GUn0MXadA8908iG0cjPeRV669WM8FFO7UPjeTfx60XpsKZncpf
Ct6bdfbbmNT79uuAbvrr9RYuxsYz9zayEw5yCxqn/rrOrlyqH4kO5oyTX13YUX0F4UCT5Gm18qDj
siEl8bC5WfF+oQVSPJyEDW3+nLadg74/jxC3BDx5xsJnsvEesAZUg0P1PVEmdKOwH7xatTgjMsME
LrRYIq5V7UqfrjKEtidlJpgb+nwjpaKw3nZAdIXWTJtWpT4mCs8dGS8FOW/ETTXzVP4b9oiUfezU
F2pvQ3J6Q5KAJE2apy6YIgZE484pGVEBxwgE70814k/Qq47oDJy9zGJa1/xOTKh3xpdPbnpEvkvC
mlFXdHN2zGB/COvEc9KMD9HZC644MUtdgBZVUr4W+3dGbBB4icwjcLpvv05O7bNiHOc4MTC/aJIe
81mS+M612GP7omtehutD5Pq5MlrCTTt2Iu0qjL1wk8MaH7sFYSkcSx8aqj9bgAGTYCBjhPzKT0MU
qTLAnkaoBftgrP1QYSls3z+EIHrTmyHIoSoPyPR3d67Ha/hvbTdFQZzsWkeWczl7CRzoo8hgPuBL
KSM3wVfAWmrkYt8xn95cv7dycIHYMGR2RiOLLZfIUTwjg49mbOr6q+uF2jBi4S7h9Jj5FQv/CHt2
C7xRKlNgD3qr1FvhzrLh0TkpkeP0ngHez9+HyyjasMSIcEucFuVGFaGa/bTU7DtODYBHOIO9+qDM
6Z8TnKH3AaFN5PwCXfUUDIKdQRIyZZZhPKNvCQnlqIdgnEQqYntO63SvTWY4RuvmjW3RZqGBAqa3
ODKEV8pYzBLPJenD8zTu1RkcMiMmIdJNLRH8JHYr+cV8Js4N+i0FcRz6rrfZERRIGcq2cARB1Znf
dClAgINIrmqRDd8SnuB5p6MIrDpiXvRDNur92XGwaK3YdHH4aAzVgZGPUR6fY/Pl6QyJ2E2cFeII
dgzUwtTi0qn/Jyic+hAqIYm7NMp1hAE9ZilLjjXc5kn7cePJTEveFIPYOpFnjCUDVS2jSrjKdLlq
6URQbCCpTZYYOBHftA4kMG3acZdG5/2IrxNXCy4O3kAWuweRjcvdPF4rYIe8DlyuRLhmdyhHalUc
+2tAmKsb4FYqUzXMtrm/e2OuIjZFqNPVFDQkAQLSeLsclkJHwWI8sdN4ShQhdC0aISAeSDpjGFN/
af7sonmJAyZwx5MBTFr8fyW6WL4sqA5LOJW3QPYA9nOW3CKMNFfZNddFNoYP4GpyJxTb4oN7yCNh
MdyCDtcE50oHkAGB0yErIsYr8I/VVVNW01Qg3kPJSzjC4yKqdroc77J58tTY3BZixrik1JM7JyFt
Q6jOG01a15a/Emt+Hxq6h8n6ZMIzs8t98GWyrOmNBJwFkxfGd76JPg59jEehgPjf4yeNkVT1mk0v
ObZDqskcXZzrOM9P5Uwu1Sr6qKZ1vccABmrVRS7/camTCE2ukjmshFSkaSKpwXpw3JRc1GBrk7Vm
t//rCZzMvGZIuNllj7MiQC8CfQhn6YAJsBTs3vBUlQDeFhIjJxr08/lTsx0Klw/TMv/t1yJ3pOwp
AdZSSkmNKArBrGJgg+wXqglfkCBH4IqSsymfhSFnHow/0uWT08vM8vAvOEwt1QljIbO0mcKbcGBl
MtBoL3fsOwy2RfV+UBzG5fM4lqK7nUAuFajKx4ddNc0qlVKnPpxwz5sCbYr/a4niMHh4bj7TTKCg
EXdBJJmVrloI5adOYvm4atTjbLQ7i+4fMJkBozzGzJlQ5gW730VYs1OztpkvywSgRe+Myg6YnHSu
EuGWtO99cMyn41lLEeMhM9cDh6kwrzil+tV0S//0B3/Zw2gK+j8IpMVJtl2sBBcPgEGZjQkwgIXA
dCiszrpJt539IX7QdR39WtAqGiJOWtdSvMU3V3bDZcStQ6mwosYUC31Jh5JxplWsVATF+JeUUeU6
DGdv9bf8A57lhvXc9EYCQZds1DyxWD8VKtCCR+0TwRXRMWIHzLAmkwt5ziOESBWSp3d4bdBxIH2t
1+5g+VX0yl4TjLcUanAY2GtA7azfYYQQm/xmW0WHkn9lDy7Txpr3mgbgwKGzZ3DtUeHQSeJOumr7
/eH4+w5UjnkDbiTdRvGKM8uZPStHMevePy+mQSaBSwo6k0qT6rc18cZdhas2WKupjfjXN68X/esQ
ETzVvTC8YArUOCBcEopqViK5K7SeY/tUwEQFIV4a3HaGdfiZkkmUQEDm2MkEqItE5coQv1IAZrOo
3zbEFMAl4JGSqAcitZ3ImHY82V0kXtx0WO322H7ZNd4rUQoSXcZlCBuUGAnz6UDZjQnuxIG/cusP
l9SyfqqLZk852s/arKhsRV5sM4qx9UuPPJ+BlosA2FNaA0NxxeTtouHc2l1CymxYmns2qkuxjxEA
1oY2pULyVWuQ8dVsGJVy3CtKjcgTs8aDO9I8uTEktOTCs+CCb7cZxutNuPZWwZjokfdQ1CP2X181
COgxtzOXA6zzoxEmTwrEi2RuPofsxnrHbtH5AV6KVs0R4su7t/jOW9XB7DJM1Yt6wnnYSnD2vyj3
CveQLFgqjzfTZt5Y775p47CvmE9w8GD9ryfetyUKUsCE5mPWR3EN4hkiXnqCAvwaqKhGsiD2ySMv
GgcMEBM7XRqScCwtq937X10j+/y/HmFClZDhfl3L+PeoxHSDhFaw0zdPLcGuRERMNYqE53sJj0fr
9EKcUV4u1YY5LhHr8Qqdjfu3eqi5cOWZmW35iunxj/P42AVFUyUCn7eSlyJ22quV3F4iGEkPTV1u
VGFcHgt1H1Ib5Rc8Z3hGkX2tum5Pj8P8jDUbkVLGZ41EFB7kGMu3hyyzT4or+NKuYmDCBj8ZB9+t
M7oY0AIHZjugsAXjhbg9VTc4GhgrraLfhXP7oWtGKKTkQU+eY9C3UlzGmIWQYBi629q0gKVflB2j
zwUFb70yPoO9pBEvXc/xx7mkIpSBvg4UWfdjqcrRQcvOU/F0YTVhQ/HwVwCzp6PDpCxxJxF41Q/M
Kxe1xUAsnZ5LOLqeGvm51utay0novlQnTZsAHcEs5jfEql/BCMJqA3jqO5VvkZMHjB702fI2bfGV
qL+okyxRqG8pqVqyPoQfXvLZFFmXpstPhqsoDNFGgh61r3duxyKqUbmhera8wmCy4FeafNWIfdjr
xl7+A5j2HhWoGSrGPKgWGnQhvjSaVd4gtORTXeH1qSXWF37bZu4XhkJ8ARHR8ozx+bSU58mxDgXs
bg9nzLaB9kB5k859gj2+Dx3hra3IX/MjUdDYqzOXSGsRaSrQt+kejngCTbWPQh2t9jWlmSaXoUi5
zX6D0TuSK4Adn2jgp+FjxGmpGH9fl0wFTrGqzWDepAhudD4n5KUhcKbmy/unNHNGixArPrvRtjVE
uRE3SrCoKNRSBGIwhUM9WpUmuSh3Ll87/WBrgOFNLMVViAX4H0u6L6GxAz3wuT/oAb90trG9b91D
vAfTJyMVTRiAyXBcweAedojJ2DCyRr4SSjrQCBVPhseYsVBUFUcjSlJHwdma7fTWv+sBLSUDfn3U
IlX7a0CrckTbyo6r2DpGSPsSaH+EpKC1cn2OLWDFnrcV2N02RVDA64jZ35OwYrgqjTYaDh280hfh
47ZEag1yo1K0v7DR9WcxNDdyZFVjOU8HUUMtlFNZxOxx+H7Zi39nmI278wwALkM2NPoBFzqiRNnp
6C/dwYwT+TUzTwInHMsav/LZx9IjsPHsdPVSMkefhnKZ1H3rW4Rrvr+L6hg8lphfbFgh0P49bwpL
Sa0PNE7r+ygaBr4nJhjDMhgQD6r1Z7Ovz0icD+4bXoEiaJSxr2Ke7P9Tn86yStU4wdONvp+GOS2u
8PNvWrqFnrHJG/ZQ+RXYeCGjyHExFTaX7QzdsaTkuGybU+XdnDnrYxM46eUvfUZl+MWKvAqfJKsr
9XfNCmTk2HkQHxwC0+bzUVjjX7lxtmKXOi3ZoQ6RCW48ZlWRA9rZJW+R3g4sArJnsyq6FwIc9yVd
dLIYcFyxx7DDK2NrEYi1Fj2lzNTdWTGlIThpJvE37QFY+YMfwc3biZqFGX0moD7k2lxS2rJ8Yhc1
DX0zJESSOhu8UbGhypqTB7tf7beTMTEA4H+0mxta3HIXDRuIT2oRxMtuYMUtitlbucfZO0S2YaRk
7t+5oDTSKSG2eFRgL5uzNmWZ7QyIcMklGLVX9CyVXicLKgGUizlgdFO0L9LH65xEcNsAy17Dtwcb
EXeJIW01yLLgxH/m99yCMSOUqKjHerKecaCBImkkUlyudNSbeQxlBJfBlMvwF73sQfQbT0aKK9Dr
K/Gr2ZoeRmqH/LhGAkGdSUkzlgVrqmjSWH7c+KLOcDCp5dYiPru0agoOK9bfYcmzEcyWBSD2ATM2
UZqEOF1xYQ+hoZQdWq4WOmFBexb302XxUEt1mw9eevtZQNfebNCpT2UKfSLC+yn6YAI7wI7lS/Q1
QMZIm1i4c/2QOoM4Z7RsPnP3c4lKRTmb0xGEXbinA0PAx6coiArRnvJ9u7I/eqnLQ4FfQK7ASKjo
8BwZWOC4oyEQt9ANhsAuOFfW75LUgqtvwEfktx+FZxYWQ4UezVotrezqv+d8sV3ETxJLhU0tvcRj
pZzXa/TdLSAdjGUhj97vk87+2BK/sO2QiUifF/7CtRTfMXxd03H3fulPVhVAuRJG1i+a79q3fIDy
x5aehlv7gcyV5Ox5D/x4jvBQ3ZYvF9sFfc4PW7KdsMRZu4sP58G+l4yv91WZREH59VvSoGcPxqnC
vEUsSU9BjHkJS/OCbbIlYHJ/3laL01f6244C8vuqDm91EyXM6WMyWJv+8FvbwEuQotssLvgX6L9E
uTOxDNeY5jab8hBefZUz47Ls/vBRwu597zRlRuxY1uqvxhZOWiFh3BF6IfEDnSYupr+hGF0KzEt0
V2IsgZW/0jwzvNQRY8THxmha3BYhIm/rttoGdUvW8isNe0TbkeL3SbV6H1G3Vso38UJIzMRPaDA4
GG5wEKEC33HldqLTCOFztEC6ISC2W/aiiCCY+847BRGSpeUY1JB2WBWleYBC2MAhsdx1ZUWB5aG6
TpsB4+ceb/LQO9wEl/wlXcgU3E2UUq4TifmGGCWBWPESq3ELPQj0ZDXreNAo7MZTvTPOYgtMhqpr
ihJt3e4x/wfj2uucJZzqLx48jB6Gs6wk0aN/hu2KZe/sI+FiEURrCTlXJKGVjkQwl4jSwhhHqz8W
r5JIFRqEpBc2LwyeK40b+tQLtS+9KRp4rDMeEWv81LC+K6BYzHAuwaOhzxH5Tg8sGqvKhFJPbVV+
d7MSciLWE9gs9kxFQItqHu7LlFxXaW2isIORnDtf1i5eJWCXKInKMmZd+JYpRwuLNYNW5JF6Ihxt
aCXjWRkPcoGL3tcqTYg/f8SbyXGjtTToZrkvwY5mUBUluanrqOX7yyF3ekYQul/nCXwptNSsh+th
XKKrFV/ydS6d7nRKa/w9GQuJbyGlgwUuSEtTuTYYTVBh9/RhHwxc0IA3lu7qUkpeoAiEqPqSjROu
7FmnXoHEU7OKa4nZLbYezh+12cNeDZg3szbQoJGkTaLjr5AKm6p1/PDK5cKuN6aTFTgLoHGxZng/
IioDDJ/G+LUbman6oMqrbi9IWQE0SG2kFRrflOIX6IBejyhXcYTz7jFbCqaRDIzHrIIRsxKVoG6u
jkRkjAiB0KUUTEdf8AaBG4+SDokrcTVUEtw9BHVkOIMB3pwQ3z9aRFUL84P33GRVM084obD+/hA5
StkAD7fVqB3djNHQrvN8lwtGjUM/uPwDGRs8TPJx5M95EAs++VbJIATKHkQZr44g4wm/1BX/no05
AQlhliM4snRfGoVR8EIn9yhCey8KWP/9wkPvoP7NQVtOg4WMqyZJ2YfxzYsgYun6p+dm8gHOYmPQ
Zhtr4fdhvFg6bVw36hThVGKPmcX/6VWQiqTrKs/TfnlGgHxwsauJ32t2QVHa8wdkUwySVK8PQfTR
/C27GiH79K8RpB6+Ft15Fuqb9XDTnfPTHYSzxSRaNSx52uGn0M0Plls4T3JxTlv5HVlv582yQ5es
eDMMlIsAvClugzfv0yrDkJt9z4sU3Qhz6uqe41n7J4b/k0oGN+Rs7DsfhTSAVLKcXRdac2Luk/jC
EQtIPtG+kx+oOI/kp/GO1TIw0zWuxJ4bAuv1EbBXCOGVFAMQdVGgqRyEEJmUYfLaLrXAVRFMdhiB
dlTCYKmhXs6g05mykq/0JstniGta+c7q5pB+qKJ+tOoOuyCTtPphARIdH0yXT5hVvDtuVRgVWxbm
3hEXOIf2AM+Z684XzXHakfnNgwvoXuGLf/Xs0L2Yswktio0mM5yrJdDWONJFtS+DiipkjPuBZV2l
E+b8a2frCcdmNv5B7HX8kzMmNgD/BNaEoSXYSI05WoBkG4VUlwzLH8tBb6L+svneK40gMut1Wwhq
RciIOc3nWAUPX3SPoaFUg8slYHlRkJ+98++6IHtUa9pT9iQGYsfAy7CwwZw+hPRsevngcNU9VtEm
JaW+NjCHW57amOgXMgoCtzqsqhu29OIBMVgm8IS9nlvkmN3IsDm0WuRJ9EIEYBFKBFeqEldEIabY
e7tRgiQeKtEgB/q0QNiKH6Pk7EPFH5dgeJoxqeWINNSjEdESgVvzVz3nG3H74DLrvoaQYH9ed5Ik
wQ0PsIkq7mA/gw5pHZb+gbfj1RtfSWwqPDBw8RsL6VWyQ/6C3ESz2sh7eTP9fN507GwRMkyN+q0x
LuqtwwVrzF8sFm2akXSHG9J3i0cRUXXP8qWM2dFVSRP78TS/Af4++9LDFFo9I8EV8HJClRRV2F/f
c1OBj/5G3BtG1UHUe2qTnyzkZzOPQS4ZNu5skS8j06wks46ScHdvDCrDZ/39sf6w1ZLJw6LclbX9
bZ8Mc0TyaoXznBRByBWfg8itvV0SAvexOyOogGGvII0R+t+1flGmv8QJFeyaSaNIxecnh43e7+3B
jxu98PupEN4rMESvYxzecPeTV0XAO3kb+lS6TYTyXmNiXfTJDhDGqxqYnrG9dEH6OGR4mUmO532T
H22Ubrepg6sDkzQE10lH4VhD6vg20/1OBJ1JXPh4Tqy0aa/Db/jVMe9JXmJAw4M1wb3wDvZXUdEm
jSGy/zHsQ34s1Goa3JDw+qEchgR1LQsPnioEEM/abb74/naPBDw+81NXY/tyTpXevnuWoBbuwUxM
p+BPo5eVLCQRB39i/8RrKqJoVV0Lfsmzq6N4ZUx99rxZoMTxJHSI2Y8tmWMt2WpJjVgoBGaIC0MD
0X11lrpvlRSRdzWx5r6LQf7jjDZxf9tBp7DovudTmRtp87m91k0fYDgHWCrRVueVBXfMJFiUu3pK
obe+H3LPTgB2UeUQp7yNZyMDYwfmAJpGpReUilVsksuFZrXX1Nr9k1b15AEgR+MaHAGmKBgHI9cj
MWUse3FU4FnbOQe0QPlxsCHOc4X/ouceUEb9ETVwTfrKmqFh7sW+t109Ncvgg5hA5/NewyOthSsa
JzX4sFjTpq5tc5I9oaPmSv1gP8HK6OPUvtjrZimlP5y19hKhYJ1M5pdg2yeXkhHAlW6v38XfWRU8
gZNOgBJrFbOgPOuQRyCj+q5V+7btr/ah0VrlH7O64f9jWjTHYTsnGqJT5x4hEGYcponWOKo5KOUw
iwvV1WnEKLx6j2xn+/puhKDFP+JEDLkTstc8hrtfzCaldqdB8o0V3wV2SL08jFgSydXTJcz7s9SN
Y82HMHOlIhSkUUVoXKLCGJTWNa/OIv5pmuvihxLkAK6HEYVilA/k5EijRcTCK4+IAN9JP2YaIo+5
Gyn2pm3sqfh4km8yhVGJAD/WRR848C8BpjBCzB9lvoKxzy24yQdstQVdjcLVa9ZvNJ30P1n2YcFD
/E1kbNeroXPlbAxm67IcYeYnX93vGWZqRTa3tHg+OQ5zltmE75aHOfWRn0oETKjMl9ZSQtJ54qBA
2nEWZKzjFiSCjpZHS+dt/xq1398cvePUjhNxRCTzBPKUPmN0nBVJDykbo3awThmZa+181WPx41Pd
uT3wr6turXy0PnXmT1QIV6vKfMUOxdzwsWeD5BBmREBLz56oyJzInha4ouDxLK0HF8SVXWrf0N4G
blxIscArEv4UFxkNxyzJKVJmqc40zHVbDVZZgAhSz/dpv8psipBJL4MPnpNCjkbise2VrOhstbto
xKjRzjy32HAYIredkTy8wT/H/1xH3YTUi9fAjUmf/QWuvhmma7GN/CWddoHk/Rwk69hIF1alDXBg
inHE5P5gLdohpROkPVMfsEx1DpfckYb5rJuZFBZf9xZek5tzZJ0R85os8cQSqjyBJ4MjYmQ9Z3BC
NOVCG5YOeOfqKgZrkjQg+Mxk6PQQaIc8B7ow2FrunecMIVTgxXJQOPp+IxISJ7mgaLjb0FWXiAdD
gPTaP+dKv5zResbTnwQhU1PdKOMMI6izg4ZDktyfpgl3uu61x+46/dOsc5rLARGg06RgE0xNyJ0r
I+wVS958WKNS/D9hYa772R4TgbujVZrWWryunnrahcKHpX9+EqZaCrT0ez3bEXoGz/IsnVdAK8VD
H4FjDt3zuzxOKh8MP6pdxhAN8xa4xkTdlvdsCwSfp3esC8jn0DQn3cF2i6y7Jlh4wYdPrLWTwPEz
FSoEUP+ckDd5ejOIjqLvVO76NymHzD1XbQjVJ3wwINS5XdwphtV4gqojW16ShGCfL08QCF76a5U3
UclLf7JyfC/CZ2e5oWknp/WS+hx7p6y1Q7JFmk2wCvpgORSAT8DOyU3Bhl/piuILDwoEpnxK+HyZ
n3ScPTjYnZ7CJ2+KuWg9iMbv4vVBqPPnvY02ptQQEGe0JiCe2NhQmGNYX60TqWOQN2HmpDlq187m
SpFwVCVGEQDCd7Y4kcqC0Go8kNZGkRssZOUGlzhwGzdfcOqh/x57LAkCaswd8TTy/sQ6sm+5IxYt
KcazDV0AXI8wMfU9sXLGZ2AwQVeMFpQq+NgOQqmFaoS6+cpAnx/BZUtoIF8ECZTcwRTRudp/+TaC
EdNtL/2OZHpjLU80IOltU7NPQ7Xu5Fe59C8uGd+HTHhuXzn6LtdBOtwlqUajLk7IZ0eUnFTW1PcE
KpU4UEJfNEg3yCOXnx5g7Q+KFo3Sh60EYARmv25T5ksnr2ZVuGtwn02GddN0SYl9JaKTQga5d/S6
4ZBDYbJ6R6P+azc0roJnuO4rhvJnwfXyt3VHRk6IrgWnvkbaVRpZDk3TPsi41wqoevPkf/E6JGOE
0UAPDfDSR2MFKOakv4Qm8NfcbyfnHBt0OkV7QNB4si7ywh7ssHWJ8Ar7wTqeGaBi6kP9nt7myDER
lzASrq/QUnTz6UIuApRI+CYCjOVf1EwxBnEVjaqoJZ8wGVW75DFh3Wf57Vsc6SjOg9TY37RNlD9m
6jKXLcCz3/lV3IKI9yqPKceAQ9AonzQZQg+HRScZO2bxX0b3TudGWppqXHhi8wmpHxMvnH49DWPA
M3qIFhWM0rwWN3tDVHZu+StUM7rmAf/dntkN37m4bgf6k2mTxCRoKC1I+FE9Ld/su5Q/hLhbGo6n
UY4Ia7PuZdd0HJ6z78ACqfn33N3bmJVLBi7ZE5sDYf4VZeTEcEE11Iv3mp1mRIn0NaeXaKVzyQ5D
brI1J5+QMRiLpXG5zVFrDNfKMyoawkuAQDxaW7/vcB32FIvHRY1+6k7Y95RlwEDUb7b0LocLRvzw
b8jiW1iQwsyxIzw8cAVmy8JKemFv6sYf0pYLZWmoqXV77wjK0agApFYA9c5mbn9Oq35/B/cTgsr0
+qW2yIw2OxkKP3tp1f5r29nwP+x9TqafDYWaqRDuVdn9nLr0pl2vt0l5ljW8JFzD7rVqMIEyY06J
cQviBn0Sw1iXrTJEY6UHMlp9WLejEpKDb4dftqS8oJj4SSrPmj8pntpz0Ftj5hH30qPIKgOq7aqQ
8Xqf4svPVoMZGdEhUOVuHxS17UWxQZeU03xoVRxcz7BzR3SZ03yGibBRsJnC1uiE6gEfQWTZZ6aR
4TYx4DHtF+zF0q4CaoozB8y81QRYmzMU9sG0uxSLLvdmiQTd1MUmJJd+YRjNlxlwI6q+0rx4QJcb
1mM6tkt649Z3fq/QBQgbn6Eh4Pk7PDuWkJatEMMq2veIUYaaGzZpHjaoBdN6Hv+ZrVRcyjXRq6hG
0jGOPmN7bRbuuyqst6LnrKviPom7y8Bgh/QVuBCB+rW3FZ51n8r+/OMdWUfXrZbVHH67YqFAh8OF
FsHDK4KBYWSsAnXGFQZZeoGISbBoWBkczzfhhP4srCA580snc6GMZW/34QVaLjdd/OeDrDOxwswS
5DiNq5w3YZjFpjH+HUsCgStB10tZ5bP7uQPsxHy8mUFLEsmg0VvzLn/OaKxGAM6gsBwW/vJlh7d3
J5sdAS8e7NBpNYz5MOGT/n87A5CKbH76bmIXDEzTa3tJkth1oBegmwgX3kmYvhHmzafX2CcgMDxA
ELr4iBQmdJzZfX55N86sJCwyNQi5ROJ+kdPjDso7UTfoSeDcEmyoYM5FLNECZtfzcnoGj3fBOqDB
BV3D72HuNnTrRrONQBYRZyjzUcE30A4WH8ZVTrF8SnhDYr5sUT1ErqA4554qc3ry0vsTRC7NETDG
ntS7xu0ZWOSCvsrkHLh7my500pnpiKSIlY9sEkOapzwi2HTWVlSBRnQI2wDmtM/bXh/Eznd55q88
ZDffIcEsDwipee58wW2kGRzWmqeGvwD2KvwqbjhbSPmAzsNL/DO4P9UP+NZeSRT55vfCKu4Vn8Ng
27sFxFt3vm4HUgxbklHIaKZIkPiddwIYyiz4Wmp9G2+lN1kCvwMiBNj9y676UFfGqQ09OE8QX9Ws
SZjDKZ+/QKYcs7VKplqdIqlcyRV6eOQV7jeA/WRWcrUZJKok9vdkJ7isKlnULfS9LU63a/UPPdKX
YMv564CN9STQ5tc4Kdg6PelVpUux4DfMfnAjos4PkERh5wJ+IycmlVzGYViRUqaSRP6vQlvDRxk3
xkddKOeYRTpa48EuRopMGfUQnrgbWjXt+HxVFjHfWCnB+iq0KmSqr1wSVM6ZL5dW0DI/T/rQNPZW
1WdtgJUa+z3uDCrbFDwUORyWxDZwkah/Sqp5uY6ft/wW1OVSkaLs2j6XxhitGlAPC6HDII9lVbeP
KmM6CCaLO+vOtCS5ntjtG5e6mEdePFxvmD2XQsDPBqMJxjEMezib5CNKsVfKJQlksdQ/m2UisS48
kjIBxcO1hGaBDnpbZBFeBKmnofMG8asbaa1DkZYtjGBY8MPhonsZXM948aDoPwNSvq6NmpexKg41
fn21tJXGoN7PfKaOOsRfN7Gz8pu5bveoENvEwPkO/9/D0934tr3UrYbPSib8OzkWMFrcnTQkFzsP
cK2JIou/xol0d0dkMRK8keMl7yuDsB12m9/vvPZTty8V2jMlDZsit2QholqbeGyUGUMF5wnL0nPQ
dGLkqCpG7o0DGtQMzUPAJ/4LYSReABMIEMYSCoy+xYXcJmDxaKLtxHEEgwH/CclfWWvNU6ku+DDw
K+L8/iClGiuQ1wyGzjSJZtaSrY2JrDjV7BQ98ab2ZZNf9i2txVb3ECE3ZUBNfAmqLsD29+94KVZs
m7lEuE1iZ67MMpJdKMdwTrVqt2kO0RNuaELpHj5SFDsbjZdGRTjUkIxCm/pzvMhPEOD0+uwFHfwc
ygaZ8l2sEEwxh3aeZRTOSknov17PgD7n1sfueW5dt3eHK5/+eEefT2Gx/tthDzkNlSUmOsJ+Xhsd
/cbtKojuoTm0VrTC7eWAUeZnTuRbxYrOPon/RqUgskbrWMzO0vVoAao+nbHYInnw7y2vp6Ybd+aG
SDGH8oUcvrKdl9FojM7Isddlz5BNX9tgqvbUVZGWKRJE0pTyZGn3JLKKk9ladthaFJOuZlt1QkeS
jQlEK6aurFX4OjgrXL1KxBwlal8FMWbvXojVc6hIXQ8v41JtBJw4NDwf/gGdSBF7W/rcyqquHrOL
fJBDDxXlB84PHyil4rM1NHj28aOOR3QzANrnFjcAwF8WCeqATo9EncmUO4nqP4fbLz7mp9mIjX4B
TumSSssPvB/vMSA7m5JguS4DixhCt1kCHi6eOC/6Y7ShqJb+NeIRNogEaVdEoJoXbE+4JGAvK+8w
iGI2SHYhLBil+55VNjnJRYLE9mk054TEZKfgJqfBvL4jAuTYArXksbZ7XbF7LoRT64fAISgMnZxQ
6IFLgU9fO+J6Th78qLZB7FkLJ7f06jeWy0BbIyYChwUo8wwheF9lzzp0YcUPn/tIzq0xmwPuogNz
ZePVY54d0adg3yRGWweP0QU2rNyCJE3HSocHj2ugkr9vkDf9aRlOZQrP0rFehYJij74zC2Rt9YJ+
hJftdPKbZScjb5HxX3ERCiy/xgFgHUs6GVMcFlAePf3zMiWdmPdTgIXpHjcJO/Tz3UzsdsneFv0c
zvJeH4ltNYJcQ+tkDYTHtxadMqq8NsdJ+Ks9yjtBdai/w4dx1J4dzy4+3xDW8pRCwcNLZnvkpCXY
XzvuYuwYvmi8kIQFljn9zo/TUHDphAZtb/Y8ie6V9n7wZzR1D+7Rm668nCYrT8CFJQSVCwN+lleL
scCGADwdGX6BRhXoP2LU9YndMd+T3ETuJGZWfdByNOYkJoEXXoSzaGIDoMs6t93sUuytHSKQoawz
6ReLuRvePDYw7IqTtTk+CQ1ecqqRKvVK4NaSNCfmnXCuTRDhdKQWXGZs5LuRdTG/DqrJM2vYlOlg
/sVmWoE3RgjZ20yttr8lF1+PiIpB56NwRF7AAXswSf2+MKRSalaf/R/HkDF598WhFN8+1Eg8G01h
cCK1K2TQeWViU9DtlK6ZpxUeTOQxr7s2ZfxaXRgK1J/Mb0IjNUQiO1/Ax/vSVYIu6kzsIM7LvFJ6
JuDEz8xjiZl1QWXUXdVU2FH/5P68ISN6xQdzz/BXkwxZukX4UJD2to8yAatX1qwTOLURiwzQo+Ex
a4DbaavdDHejXapIW0gZVBcvaQs3roskuD+2gtCmCOEfb8LL9LJmiWjevpbGm2pMRmU8KWHkM96p
FhXrshXvnApSJs5+QJvBFn7st8pAzM4UYtXupH+KqGQBwyATiKggHQVcJDUf/aFaA6TQ+Bi4ql44
MhU0KMI27RjkcUsIri3lu/9Kx3KD/5cha7j6DOQ19VYqcmwxbFfX8jJg3phU/AliOTGgDHObO2Xa
PvsWNG3/DcHudDLkT0n/2YAUtD+ZQheFEqn/UM/8ZLCnhNS9ERaSNg76e203EfqO/AcxdG8Wb3Ok
cuSTerR/5a9woVEI2YKCD9uOkfD1InY4HA931cZk1Q5V2tbqMFwOX+tG1QmgnAj6RI3nBYPez7kw
YKOdCBlg0k1D5NFnlClTJ8u1Zpc6W4iiiTU9n6TZtj+E14RY95z4xq9OPtuVvyrA3fdYZ5t3UQw5
eoiMf7XTr5Sdgnq/jrx9xzIUxAtgdlcLVn9V7H/g9UIJMRlp1ETYslY7P5onfsZvgiPFP1ckczjw
TWqUwMAKMTwVBEiDH7d7QkNWEFCK4CvAfCgxC7q3pIJI4CpZhthpWwm99aDcB7kAQXqvCysMrM/t
Ufb/Jyqe9Vke6pbPkK0K8ogMCjgKQi20YKxFRcl/Us1v76vLn2VPhum1JichLG1gLI+6hArqE3oA
Y7u8AbKuUk2802VpwEemsH2szDKNzvuVXXUqq4Oz5XTCLvbEI3lYWoSwIRF/xatj9UWXx5mSf0HI
xgI8v3Yy0sRbsxAcb0RFQg0tiON4hRmq4ytJeIY7u/TlbyJ2hjPdLHSllRRgxt3JWMS552CAfOJV
qYI66o46mgACafYqv3BK+CgGgQzq2AhK1TFAb1pbjSdFQsSAn+hzb0qel+3l4AuRLqf8pQWPgyS7
H8eiw3LX703z/W3NbkOuYe91toONH1l1B+vn3i1HgsArIVLLhkkJyscnStRuGKTr9rcLVCZLvxHI
Kz2eSf/Jw6gxQ6UJFTPXbHskjDvCCAZpcaaW/yLm3xqZQvoK9vTjm+gzCvQYaDJmS2geZxhXzcET
h+Rr7DB2pNsyuKJjtEG1HmingMV7iT3a7tZ/cFb5xa/jLfsKvVGI8gvzp9dUZKhkaWoR7A4+vmvH
qCekCCV4iGhR2JykpqjMQei6i1koEbVmINjhX4bc9iOkH2fo7NmeqNWlG1qu5g1Vsg0bXiTRyclz
TNFoNo5qFQMw9MQxgqVpHt3Jap+SOJPuNzaQThHYZ18i12fUjVdwtYZiNbCxzDx2w4f4V7t2nB68
ExlkJo0yCcHvKH+uay0HagGaKtFRomFeekjVwAqGDRER2SuVXiH/4VGliXg6Y31DN96ZudtJxiLS
Q7J3z2HUimydptgB8uR01Ted88hK8hhLKsL5/57p2DgWMs2WvIvMSXcH1+LQ7p/Rsw4MJLZvNstQ
72rfiBE/0GKs3xCMjQEr/SufupD68+15YauCW4JID1rBMeiLJiIEe9BqXnI5+wlcOvix7Vqm9lBZ
G9EqQhx22hYp6JwtsJZe7xUhdbqBnESWGrxzGsFNa5QuCAkEB7KwRA4oijCGD1DrxA2D8sJShPKN
S+wWqGSvm8RyT29NNUpQrp4tgJ7gizHmykTbfjdp1tt1uhvv+EDSJ+TosdMVXdc1FhN6QjGgCNfA
bxgS+u65dH3fze+geepW+uta75o7LiebO9gLpfzrdQX5HsgpP52QAh0/ZoivA3rJYyP5/OUm7qdl
Ive2F5III067q6inhLayba4jsV8iaCQij3VOV3aMGlswwoGDJJJPv1HYLnPYEzu0/5gFgZyx9KM3
7XJtuQaNKisK8Ltp99TE33KMXDNuQ7yXXO6JumKNP0fIc7rKaImeYHedjJUNvnMDhcaaBNMElsYX
1OB3+DZNibRvIWSOVwS49OHqsbLEFEX1JkVOTTaMoX0QUP4kdL87wkinyMQmzD9jMtI5erQslYKS
KAzirEypknvZ1hIyZx6n3fxouD9VgCWFBHk9O066O6E/Ax+K+K6x+2XeBErJh0HD8rVwuRLvRECW
LjzIKW/Q3MqHUbeay5fttX6jUO6Siuypa9yGJV54JIXY44mqP2jlxnCmjCMMrAYnCfM041mYqWm8
L1xQQi0zd9raIlFd72zEq+vwoNlWVeCYNLO3WgViPYLMbEjtaF/8iSFfo17iJSIRDFRH5Zlj3Ypy
j+TJXoI8NpnJSYdnelDFZA9/osICo4bDQCgbyhexoDEVhu38Um2LYG/Ld0bwHYdwdskzgSlqtGpX
LiUikIeYwehalNRQEl+/Am6v8o/YQgY5yPKfqNCYksYHYOqF9ZzYnXRshWRceC4NNxqBxdzTRzlE
4h0rFTpLmXuW66Oy2O5QqgrLMIhmvGYv2lqA5XFra4sOHs5pfcNa9XUBr1ZNq7ZWWnoTphOhF/dj
eUyrR8I7aGCVT9YGR6i9XLx/OuaRQGYiuleGTK3jjroDWat74QnVYSKPWnPWmW+u4bGiTsq6PeYX
e/yvOrux5r2Om711jfVnRLyDT+OK+e0BeCQMnXhXChxa/F30YCaA6eDYkDMh/CmkUJ+hHtY0DNL+
Z/yM0RQX627KCN6UiRXMGJNt6X3DGQbiio+1giniqfJyZ0tfKfJJtS1criAw8xP8PbvgEApg50pL
zVVInEsmgqLplu/XD07UKEU9n1Cju4fRdcC3vHEuGs/iyOXz0zQIAVVJnmkBlu1CZTB5X3VDX0S/
/rilr96VDb7G91akat73vc4GG0v0a3upsWaL0si7LBeIaFBlNeqgUsARiYFwqub9s1o5Kfkvnho5
1zBwquZFmPKJ86v8Nku6aCnFWrwA54GwfCZ+fmfCizTA6P7//s1jyU63qv3J/wLlS6MMEQ9YIk/E
yZ6R8EE1fewNMxrya3i65mNWNMXqeCJf59ab+UycTdUqVsJAJwC77xrAH1Lr8IHooia102H+FB3G
w+UJznx1S/Px0NYbQT+okQd8CwvbbUObDHfK/MiTGSLY0NIPi0RTKZqpHr9k9LVSNMXyB80A49nQ
LtsX2MmjE6l2kB4XNlm2WmSCipOcjg/tMkYv5gEEk+xSwfV5mk7qj7vbhAVQTS6ha7MD28DSQV6M
L/3vu012fo2fDDtpKyH0ABaMp9Xbady/8a6p/jbzKCvv4vaZl6ymECQgPKhfLgjykapYU+7TrE8K
/5zZF710qJyL4le1nzEBSKH2oX+LW9Z1lTvMRvFweJqqxB1dqJZwXmeq2i+vKO8bnXsLpMlB3qMv
62gJyJR2MnH7jM33sr9YMneyhDIfKhnhipKc0F01+RmLDbNJwQYVI3YbtNY6qfZuk0cvQffCwfAs
pUMVpwOu6ITGPTFPQ6Ea7nW2Xis2WtjSHFXRWr0XooEANBp4l4NuEyaGau9rOgCNpLNOvN9cvSyw
LP+furBzk1JNizC0dlmJh8DtwE8vRqNiqtmzaMF6OAKnWwjzKe+siwGyfiDt7S5qk+qSTYEALxEo
9Iz9cEbE2m2/LyigPSIE4A/R4dOJoaGBPSy4dE8W2NwJKpjPlwQV9CIyzO4JUQjAmg3JLa98D7I2
/PlE/UurUw8G6gwS+aZ5ZvshHw88DZkpl82YZQXgMPIXSrOerCKhLDO/wcCD1GR01YuH1NT3R7Kc
8KJwf49nMyhTrhjgbAKgehzCenHhe7GPOPh9UHIA+vvJzs2Sq1NRqgSBUi+UIMCWE4WIsgnBrcau
3aFkQky4xiPhHJtdjS9LcmgCg9MJJimb2uoJ/3YaLdEA7jlIJiQfEcXxrC0VW2QumV/W0ePjlLJw
MLkigripB4YUdM3FzWm2r5mWvJBGe2KXQoJecEQKRIStRwwyUk2uxLQMM0v9OKKrz2ayxFTSkOMn
NvTVsbKD2kOdG7pffKqPp7grj9C0FxviLCOFRrrvz5DhoqBq7yg+X7spjmaptPKTud/2KrXEZtdC
RY5HmjGJwyZ50ndFeWZs7lppL6pM5bNYxnTcxWiuEJYdOGBAtL+FRGhCj3S4UgiyGU5iw/jrZR6Z
9uD6q+7cn09SAQ1algUpK1G8cpnlRCPdYvQRuVwH3nusYhdZ0O3eYs02RY0oRgl5ErZfK8YZ+Cwl
nC7cfN1856bjhv4B2DPN6t06rQbiVj5dp4Q7u+NxHncMBsRu0fjrxIHLb0SytIzaZWo8eOpoDPmT
WCYL/NIVGRx9e5EPxEav7SQt/zpBqErRTMrk6Vsnhn4p0pN975KXCgNq+OM6LUZyNMKyl1IWT2Ye
YCb0GyPTIARsDZwmtnlrs5UKPEc5pHTf06gKvVU50cCuTR7IvZPlCfQMq+2FME11umkQewQFRnrY
izlo48tY2Raax2cKThwXJ1BE+nGkT8X71bo0MDav/mefp9NJqbSqu5pXUzC0fEaVIlVuNuZEmafI
zK/Je+7rrVfA2GFbyH3CVGIcaxaBaebaE2pY4Ct+lZombnAyfRsJ6VlVj7QCNwuGo8tX7RY60k9+
vodfXDi6Jtp5ZUwnt6lB59XGiZeVGwDj7doFBv4sWKgL3B6amLgb16g4zyeoDY5aYoJlEwrnT9an
/s0p2t/hmpgGoz/ECJrv0zd27kCwOrrKweok2kdrfGBu3DMel0TNTDSx7ISLlZX9jbyh+Fw37piH
+q7t15ISWZFWF8hwJUm/g74b6BCcUDf3WbMqSFT7hcaM8tZ58ViLsIxupZG9PTw8dzS8cE4NqCZI
XW6i7pa9ltCluIC6IMc1BFCaMus0lMsNPHmSZD66IeTge6dGwpWEy/lgkeHYc+2vbqZhdLusoU2H
SJtXa6kL7Nk660mwRmsmj6oTTObdMyxJQgJScRyKnZ6z5VJfGg+cmAgVh5rbZCC0DK3lBPeX7SNG
LL4P1MOdrbfcFfeZ/ZbU9DzvM+MTPlPohRZz8+4QBw5FkjPUiSLM8O13YhFXYnNn2jRbI19N6H/b
O6TBzrPiTBkjZA9VOrQ31l6zmKdVhzKy7ktS7cbRyKfvpL9X8F/ZnkmKD1ExA+oG2sCQ0V1uYopi
pgMxz2p936skTw9PO4WhKiUh3lKw6g6jV+b4VDfoJpriNQERvw1w8R41lapp/ROWi6he+41lJDq6
MfWPNjcX3Qxcyg3O7c5pYTsCP5SSkr9X912V89h2siQuR80Q6FScr8XFgfkCIH72WKOeo1n4yBSV
/C2UyxEzS4HIL/pCyEu40N3Ld7CgTdxQVHOuGx+AShJ6FDkW9qt90Ho4AgYrJ8GgofCIhwF42c1x
NY7s/WLQerJJiiowpdN5zAXTBnFFgI0sRHsdsPrQLcFWtfB9mUlmGl6UB1Sz79SDK7YLIOZ+E3oE
QBb2XcWwNxsJVzZ8qa16HGCXk7pttlbnakqusKmp4NRgEqPghZ2261LeOJ+k/HhADqhy2w+Etjlp
XdYokR0kTjVztf3j1xC0RvqngISk15fBcEYzBi1gbJVex5gpagZnvfFA0brPQb2NsDNMa75X/2Cw
mSdrYibjxAbVJ7nEGeIb1RyrPj7DEi6NYI6J3rlpFOkQcxIj/TZ5nLHkuYwVXUpMPi0GhFpq6vVv
dzzP+uZW6RtGw2iiPgDnRUNC5vDXrDcxG5ULiE9TPIDrQWYJVZK7/+MNhDNGbaamkQ4wt1v7pkj2
o62QoMR6dgjfmF0ZVZewFoBaBP8Hvlw4Y0PHgT54ydh/SQS5P2RYIxmfKY7xIsGZaUzKrc5Gp5ZI
yNdEBRyT0AtN2h9sev9X3fds8bxGctzA/SPufptu8kZ4TyCiuMOgj4zUkNVa84uA3Q2e1FvHRvhR
oRwMo1mIqqKkmCGGSeVcSf064UDyM4DuwJlKSVY4MlFLoC/sbCyXjpgqc0PlKgI5XBigbBgVwfds
zVhjIsUd7XrYUUyz2hmMRExivsfnM9Vn0oVMwZmyzpFIbS3PGSq9/qnJhVAKbpTMl/8m04NAzKLb
TchLZOLm865CTfQm20GC9n82QKvkjnX7I8Oyyp5ib7l/ZAYPMzq8MkJNsAbpibXapYuixWju2HaA
nd2l87HE5s96vlg6ODOQHZCVupJmwUnxCUhaMJxwo1zeC+9XPQH2asjyVjIyDDArYGbh3q9Lx8QK
zr9CJqBSFduQ6hgUQ9zZw2+jlP/qI/jjlv9PEv5WMB8vNAwTc2dfbvE2KAuoefJ1MUfpQZYE8TNX
w2++eSIZnU2boJ4bakjIQ/wM+ZPhT6omDgfmN+F5wnZh66mfDmtYpcJ5WjpqDfKQuGhtqMlUGLdV
UCfe7TAx0cnWqYm7vg/CSuftqFAnQTkTVRjU++S93YoMSmvskjTNlC1o2u+nK9TXYVg83n+y+9a5
LXbxK8InKTni4Q4Y7tietjIm97F2intU0xYCISFXA9v/oqqn5t6vhPj0DAZyOhBAEomFfrkaewxA
R/mfxztO+lUbITVr6LFmxkKCMP0JV1bw21Jai5de/QJ/cdpX2vzGH4PnyYNPtMa0X+JUmPLmy/1e
wTaharFdSXbMdGr1QzPmvMS3nob3VFh+jcjs1Uw7GmSmXww1BDeCqozUIoC3SZ3oGf2HYb/VmOzK
SpabZ87KUCHt5WCacz6JA2z41I9JGt6pWz3Sh+fgKb+7r+xr+9Qxsy5mqvAjsUN4HJgyZbxxV4w0
A2V+a3xJcVkvy9fjBIjwcxI63Gb1nU/HiQB+Wtn+RcBDQUbw9yuvc+lfAXDT7YWV6z+h807vZF26
IGcJ0h9hXorebHjZJ0/mJyOdvZh3qVCohjCZWH5JNnf8MwMVkXTyzK2XMgObt69KoTQHyGCU3XkT
ZPpAkddnq+XPxRbEGaXywAdq3kV944hp86wc0e1NvdjYTmnppuyxT1SHZRmdSjEhTZcRlVoYknVm
uUiRr3ICpoqHvsWYm7YRuBjWAyhmjZgs3zi6zUzY31vRfzoP1Rl69fgHLkt5Fk1Lm58oLY8yuL7F
YV6sp9JnQDQjqqzDIWvfxEPPu5VmbNEaUxnsVdOmJ3LZSiVwhVYroxt/2E7bozbXFlzusu1WKGiX
HDgAWL2LbmPHpt6XdVN0cqGEl3Sj5bFyd0X3hqgWNMk1rEwCPXX8syL5GUt0hcKErHn8HNK6dMvr
DkjEQe3hPT3PqAsHdKhkohPipNj27CZFrM+OxZe6vmwgT/1cWXgL6gvh1ns9ST2ZIUHaKi1s2iOk
DOD+Tshu/IarDc7x+BTDiLNdPcAomc3EKlCGRPVzNAswrw3faVcntUqumVaKBajMdxmqGQ94g3zm
Qbm4oC+PMEf7PWu3+uRmLuxhpE3+6LHgXJVKZOWM7qvLrVLuNHpcyzY4OFMA8WRYRLm2kAsm0H9V
U3CtEbq6m0wWHojKkw2wSE4+O073r7zcUes+U7bsTFCaBXBfjG2cWGuhuF91XqBcM8JHAmDOxdp3
jmBVm+JWrXnGEvdt3rpFslMjfy3gprPg7jBr3Bd+5dJMtY915gV5GPfb7YxzeWX132hn8y3QZPFI
LmWCYkM7t9H5NyIbF/ZFPU/Y84nWhDFdjNxdKYeg8iy/2FigOtukAVN1WIiyV4xnmRrSiCNLl7X3
/VbzhusbmVmFT8kkT+VWlrY708jQO/KPBoeGMmhglSk1Afkdyegi7+PSW9W5fVNCS4d3uxAx2chf
aZs8GXhd3FhcFsoXQvsHwwi2XMmZpLMcz13SDhY+RCDYjYSnO+9z6oROy5rXY9KIhqdg3oCBViok
/yRjHOPOy8jebYVWLDI9MCFVS1GYz8HHuhgV2y+w3gDNGB1vrMdvW1HgAv1H6AMLXBlUlFbvrDyF
KZqP/3btlpKgtyPEyRogfXXet1vjGnsX3N4bDBWzHGuK6U3ef4AdG+pZ9nC0Ij0TFh023465WZJ5
+Otrw240AEC6L0PCk3mNsy7iQ5IqGZfe7rle5Faz4ZsK9/Ol9uMfGIdL2ztRaf11Nw0MKCVzOIlF
F4WKjk7vV5qzlIANmDSKQZHYJ+amYICz5Zl3B2JOkZLwktHpknzvIbeGx012A0r/cdzitDRqqwmr
NJxPvI03srC2AoYZVUa5K1PFjvYvPzqdor6xk4Gv0RoEOTt2CgSxhji16FnYTXx5TOGZDkG10sMO
wcABclKBlQOnSfXXawUyOKmlRH6kZA4THN8oANZ0iMLCo3/rjopc1AxoJQbIu4kluZbvijuQkLog
CHBBDJZa0j1vIMZhaat9LMU5GuFuqwalRx840X/BfLUBQs6ZHYptz6SdSzxVjMFUp0cd8g7ZWsir
0t/OdkM+ObWN8Nx8TGHSCjIbdtgNAM3lv3e/8T21BoQuE0Kkg+RZPJeZb/C+zx5SwDzMK1loTx0r
o21JZlpZKaGKsh7lh0GLpgv+ltvD1Ix+NTLFsxOXcuMJHUAg8tUE1e18UwsIFYzhsVHAWM1VZWfd
mvmjhQ8Vb9XVIS12ox2HD9Spm0V5w2kBJVqwzXzQFWZvotX33ZLIBG546GdNCxPB1CGwUe/N2yvA
oakg0auLBvWvBMjpRmv512jo0uqcpZUzp+KVEwhTk9kFLpimY/aezJFQrT2D6WgdpDeZnZNqpAJS
kDhYZvXc6MMkdwNOnntqomtNl4B7imM9Fbg4R91WHsqi9cHY9AM585vEGoyqk1TwV/KOIdn1h9Fe
gUu10FalI+iBiF7eWi1cxtBAlDlf8FLJl92SND6AbCzwNrX768MRdB/cazhXxRR/GYvEu+iKgcx0
/gT0tMMXtU39jFIDjQcvq7eiZp7jP+WhUOvxTXxvC+yUKCJQc1HTrFv9rf1jWNkSVoK+Hk+wVQLd
dMXRzFGuBhtwzrnhTcepm66FzSPoL30j+cDxiGmDhPTecSw9XuCh8zWNn03lBy6klDPdINCNKE55
F6PeA32dJs3og9ZGEAjfcLdzk0lHuuCauoNiUh2roKHzaJGZ8+w72Hdab6IFvPXbUkl+VJtGmoxg
574hox++q2RAu7s535aw20CdgtH9mnmJ8tJyf6meDgguM0xOlwqLuDu561vIY++Y7pwI4crTQkhG
nd/w0pcwVWq4xpWt92L4T52Kh6Vmsa1D6o6DlKZKDwNTxge21AW34KRocbcpqXow6EYrAbuKO6fl
D8fOeXXI3prhsMmHvaaKjHogCqTLQpSwWCLBb2NWThQm5PMCuTUT07sUmNnDuis2BfcxO4knSKWc
2YMOWHX/EOy7nEbrlDqdHIIYTYiG+UxWqAzKi3m8N7YQwwpcCllSvT4dXMPipG9aEiwyocAgEE6m
O1EXgpGE55n9iCQYfmDCOnbndX9ZCpGowAYpuVobpDz7Bor/8D9kjHz9G0/hTtVS2a+uYlr4kWMc
6RzO8BgXgvRb9qAq7l6m3lCbIzMPlA4sftGSjpn8nbuI/ZP/2iFWnwQoEtwQYa13VUVYTsjGZxsz
Sa9fN5ku8bcBM3haEGpnHt81V6Q0Si5FSk69snrp/QMaOepDmgbqvUrHYAb1x2Nj+lbEG5daoJzi
he/tlXJAI4NUtmi2u8InGJmq29kvOfGUSEqPoHxGQG0KhYa3B7k7b4vx39m5VTy1sUjtlg2/u1gf
XQk20MCOOgw06UEcIzO2uPBFAZWpearqpqZNwYueN2z46cHiYH9EfrEcq7LQjEcVg2QX3Ub9eq57
XaRzdMuZ
`pragma protect end_protected
