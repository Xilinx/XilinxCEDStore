// ////////////////////////////////////////////////////////////////////////
// Copyright (C) 2019, Xilinx Inc - All rights reserved
//
// Licensed under the Apache License, Version 2.0 (the "License"). You may
// not use this file except in compliance with the License. A copy of the
// License is located at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS, WITHOUT
// WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. See the
// License for the specific language governing permissions and limitations
// under the License.
// ////////////////////////////////////////////////////////////////////////

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
N4rI53fStxegnZTnoJo9RV4bRg91eKap1wBUsg9FzM0Jo6ledQEbubwrQY88YBl3H9+Vln85SMXm
kgEJ/RW9ZtU6kV7IA0XzO25ae+JkR4oMATfEiNZoKwz7PcrPD7kfInNcyiD7xOonKOVWxcWwNvM3
ZeUDZyLA2LEGEnrecEgWGdf6aGSB6U2TLc2gZPk8LxlPiCf4nXNpyoMFwhlfIAJOkM9KHnerB6bJ
nPiwa+olBLltG/C28b7V2vXkGAgSJGZpWKR/U8g0s6kLKNMp0Ojk2+MgRFI5MXcjSbhPXEleI/Ur
7owWeIm+cRIrj/YNwEZMCP9DnyT6//+BjS5ecg==
`pragma protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
cBh3hA9u2kER71l008TSR7BjkXhhxJ3zi4WE9VP/e4sId+Rl5iToZjbCOtJ+9j0qAU4jmTNHWM+F
x5GW4M8k0R6MbaQLkmMHW4MHyqowOy2WTrAFuHZyqp6PJxSRd6D1gGLJMpyvrwmPoa0dEEZosLfs
PCizR8xRHtcZH+3xmc6O3HUCL0Pj03kDuB74DbBAcyr91xslcs8nWWe70+7+nZzs4om77/1TNC1E
Z6jqPiXTjG2LOXt+3RYjPcjaHcooi9Q+De6OAavl2JfrBGHlZv+mIPLG0weR1rmOFQ1v28joLLB0
iOLYmqoGAl26YJlGi0w5t53lcGHEIRk3OylqaA==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
piiS8HMNnu9hDZD0GaxylpxP2MxwSkZLWTegFYAAcqV12Lacqb5C0G7e600HeY3NoxXuBk14+3ya
0EIto1FVRg==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
oUAe8K+uVb6yoifXqPfS+RKic/ErA1ZJ/lMZ1CLmfw8A66cQmA7ySNJ/yyadrgKD4UVv7V9hvJmL
7T4jL7kbgYtwPOWitM7OIZzqsMx1waEvUqYcc3RtiqHoOAdT2+KRKMjczKy/LfJYqaZEq0Bnzl9K
0D7W0kxI+rVQicc81COiWogkLRQBXdQ69w59XWUGgzmivgUy6PwYk95PB46ZabTNnk7Jh3p0k60x
MIvAm3o3svFG5ufvKYBetiUwH6W5SkuhcHLQ0yVOzueHAJfD2gCJvTTXRwaPBY/e6dD9H7G/BQOK
sZej3tRSL4ckq5EjiGpGOh/CcKWT+uCp7QfPSw==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NLCOqaOH2YyZaFn/VfoVFwad18EkHW1wtC7GUQzYIthdgRBHjyvx31zIbWf3caWJm8lGuqqnByWm
RIDZV5qQnHsEOJXSble9MHSmZqsKJByFkdRde72vnJ7M7VzKgNvc+v2RfgLRGedKY6T3BO0JYIRk
2c5CMcWKkU+qE3H0HaQ=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
E6fWCDiFlcdjjtOEJUj1FPhFNgzyriF+ZcfswLRJnJ0tA0HqdX5A/vqH7Qt2lxMuDAAtvU/XR4XH
0pzuAuH+cqmwMfQCJILbzzq4WyD7haWUkDQnU2GWrQj/QXhKz+WC1+2aIPwnCplwDKhD/Y02NhOM
ub0wigxfXf2wY9PvFUCy01b6TB1gUiywhqISX0ZzhcYmNX6wpEiHFB5QWtJlRBXzX57EO42lV8xl
LOj1/saACvEERJ7zRK2vy+8gem2DaGIu0P98TjVU9rUXBpd/P3BggPHOnX8dae3Sf04821vvqrG4
1Mprkoy0emVc2wyct95HNaUAEFG2QSF51muedg==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
r+m6V4/7W/q+8bT/EEgoBncQ1o2ybCgbCPSGL3mC7xVY/gPvo6kIkv4NszSikER0ZB2GDgy3HjlN
EGASIp4gn5Ie+ZrBidSxAM0TeDwiWQYUgsj15cZBWG0WEF5qjaDISPAkmERhn3RgsCAulqIAcVKi
7eT4okndP4XSXMW/bmtZbUK3HYF0emoZ64fBVQvTl60g/p459a54PlZwOaHOzdlgBFF3AY5pCHNN
xtTWhNJ2arbZkA+i6JQpvJx/BMZE5UXKMVmmYtLav8TL9XNqCfvrYGrPxRTf14s7kFRtZxSbXask
tawe7jzeFsQJyi+E28h9jP7+OnvgtQgEhQCkhw==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
clVXNz0nDysflA41/NZjJ/LzPMqjP5+vBvRmLfNvbcrUmLj2NgTZtZgY8ztY7iW7aJgLHElkrS02
gu4RpmY67jAFg10L8V+0LSnwvzKC+PzT7LnXbNFKJXNpzenv+wnHpN1qCgHjvtwmZhU0DbU6+iCF
u8HZPzvEPzxpmJ+c5+Q=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
qmOcpuBJaIOXoRd7r9BF2SscbRkiClqGCTzMH4GOoXbsmSrEJZEweG2WceyngLy8rZgfavXuSvIR
DH1WpSw0T5j0RsyErOvrq7iPM3r9opi75zXKGPl1CKeS5bk/0Ro3EbjLMpaxw3eCbMs82WSl28jC
rgJLuLidhbSzdIZbMxQfogANXyiGvXNmTK1GfOfnzCBfmzSqZvCqSktlxby9MGRikVtKVufKH87U
2mlc+uTkK7UdgwxH2JHvxAi8kg1P4TSGVWo2SqdKiCAwXNVUAMEWEWVWHDOYWd3J0Ex7xraIJbuT
OK+DVQyLJLI37a1pfXX0QKfc+K6QWWGpLKgk4A==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
soITYAF0E9RQFM1tiAu6hb8612CihHoFFNbKaTppF2VTxs+r2BG0lzN600INokdpU29Fup56pPv9
OGUCJs0f0s4afBXEhzSrzRNyP8uCGFu8lXiLzw9cm1BttOVEYYMyb3VmuZNFgp44KTA4PANb5DHl
0jIdTdU1enB6ZOFg0wzNFRwuow0iaFxqpBTctUr69C8T1q6mtM9+PTH8+B/Pz7j+7mdpeMFMZfsU
Q3OdP/fb+MZ7HJasv9Hd3zhifBE6xvmvSEAHYg/Lcu1MeDTj0PCfPO9OrWjaOsEC5+g4Pw6KFIpa
K54Jy1ZLI9CCJmhKa4SrvZt7GKLuSXi4NcmTrYWozKbOeNTLBQOEbjmtmUfAQIbkdU0j8rchR0/Q
gG/j7qnJiBiOY3uuuANNigx/5itbQgfO7BH3AJpm/rhjq4uBMndIBo1QX+tWpTDrtTSASbnAuqi3
Znq8prhU6h7JGCtJsX6WP/+rtNwnw+JjX88kQ5xHHeL1Yeg93Ay+Ig7r1T1/OIMk0+9nS/5CRqbK
/TR4Mz4e47mc9Gt9s5fF5o7NFTqi9BCYpqF71e9f4rCFZQaaMXCXbxrBBLQbT1RulCjRpZjhXPyj
JaQatNInzqETyz/0T1sV4fONtegK4PSVl6C8+1FMx2HNZBTfZ8bGU8AyDJxI15/iRbxJZtFiwIWL
uUCViSUc2uXIf5Zwb3E4ehLbKcxVcQ/5yqJb+c8uW1TLD+WajVQ+EF52KqV4YGlFT4u2aJPwGj1k
/Ng4mYqugTezW4lP+xOIDTyM2j/HBmr9dR0omplstKZ4IRmhi09S3nX3nYhVgftHe0L9WQSkm/MR
9W2IhhnOTwiR2Dt2SIbB7QJpdsFEVkcUPEGomoivgZgPUm3hZ1536ALFCb4gyZ4ZhaDY3QRGVdsw
Mv2+EfnBH4h2XMJ4LoCHWsNUVKnpPemJIJKeHTLCzLMVT56Fw1lo4AnRdWp+h0uRG6dMaqG6/FmD
s9qNV7hEyFapYFN9ASf8lIxTMnjtNstFeXpX5zaL7mem5P+Yw4It5JQrmU9vh0YKAbkNbfVHj3D7
9u6V3ri4AvTQ3pQc2AaEvWI3oZ2/SFj8o5BCtW5MCxR2hrS0asbNgwpg6DRWuxCT1BOIhj84ui+j
7SHQ1lLwkBh8qxScE2uKGYTiPEaJqIJy1X7mPEj81D7/4rV72APbJ+Ix4Q1Yh/DzuRfLShSV401P
shbuLQt+g9YTJEnNFRSSFmNvYdvLWaswGYgmJIyWnLdwP3HbcNxKRT3iEyqDpI5Wxv32jFCD84hx
8HI5d7qM8uY6TLKQyh3G51W1BMrfYOmeWesh2joA/X3vGmdcil0JH5QMitkl7tsyFEpQZqGHSxbG
raHW/XXIJdK/Ztw85eIqbkyqfKSD01DlB+UVqBn2JC32lqdvZIa5C7UmakmHwHbibBDAr1Q4adUT
1ysjskzodGKYOytWo7PYaMjclMaYS7VrCi80G0A4cYNpRnghPcfD/+lP4CZB6MQjHhP+utQhxMY4
adpB1WcZxydIivTim5dRh2SCDmWwv6uq5CTxNr5F1kfU9utfv7kmalXcKBl8ljcBnFCO8gefCYKj
7uxM9ugfNknDjIn/mkJAbjWrAIwZhC7fOG2pKwVygsEf8ql4EYmlNU8ylLfHaNH3IvU9IZstpVQZ
RtQDClDLx+bSukVpNQDjj7q4+nM1lz6vL8vFjQ7HOCRMOkHptaFGqZdXG2/IhsV4r9c4EjkX++Du
kHDTSOf55T04xZpy1QhwwQZ0TbxdY519S4s3ztjHw0dtscApQCJuijsFA50o8HAUo6SQWGJO3JBk
M0+jZRmmNMO7tB7L8ATaOr9MMgyFD9EyOLwqWz4CZBiTIFQAabj/+AZiAAQaTjrIWxXf1IyhYbpE
Id9TKn8Md4Xujt1qxpNLOrQiA2gYV52izcuwU8EN4Q1Owwl8ynjghnL+R8b/JKCmHR4BrlO/IRCW
QcLzVNgUsCAv6/dRghOJA6i6Xk1+3Em7zNWSMWMKFLLHVUldFRtsOxFgH/bu1BAD99TyKSlKrziM
abvPmmQynOrJ0A5htSFGxWTeKgDbO2Fh0Rk2/2S0lg7wymA+Qteq/eV251Hfq8oNi6S+CaYDpClf
+DEHvG44nBYjYH6sNyn5bPwqC1sObcncu4vD595D8j4uKtAV32MxWZG98hPfVIbVAhC91q1MzHyw
vPB7YqPUbuWIHZ929K+1octonwQMvZSZNP8rtOq8qMNJvnhQTNenOslLlyRxfgOe3oVrjMyNX/p2
Uq/Lna+uQuo9/1wIourVzL2kqlPUN57vgiiHp4I49fp86ddnf39kyG3oCiOUAbhXKqHj2pzO9Wes
4PyxKzVvRYrole3LervjcyM13vCMhUWpKsd7z7yLEFhrmk7cDcWxt8GfrBlrXj+CyjXXpJjhaWBO
o+xReUPTVX5FuVkWqzOGNokkLDrYFOTzDY+HxdOVaWoTym34lzxoKyjab663bvlxaqumvPaTvBUf
zDnm4cdExze1nZEzagPKEwHsLj07Ek5zPLeGKPSLTbpIXD/klBUYkMwc0kbAn5ILV7kJBXoA0lba
jJMB1ff0FhvF/dqE7e28dhVM3Nbo7In82mrZFe/NPLICeItYJNC9FQVbLJVA0KVEaF8HYGt2DTqg
duuxMsAYF5eWBNOBDcwHpL15DUe6PLAOg62oR7bzfPOcIRG/fVdexWoQzpPhvOsEtoYMbP41aJlR
PuMWYMKa7SuwsidH7BDNraaHdg+YpXiWEyQBUe6g3G2VNf8sPoT7jnLd9C0jwe1g6XijKMIh1kQj
tf4AQSxEEtlwdtu3/41HBYWewQlVaLjEI0xrwozC1pDyF+PNUJDbHgZVdLL2FpncrFBZ5zZVdQ/t
HNitxpZFUVKB8dd7Yduo8l8MQVuzp/hjYCycQTp/yuEuxC9KoTegZiuEq/GrhqVjuv2yM1roEakH
xPbwmwrWKBccF4Y9ccKAnLRpES95M+KW0G7XY79RLqINgpSf31v86YjHtIAIRwn1wJ1Imrq3KHIn
ZfHBP35mqNf6YuhzccwCvp/oNOX6c/0D1lryPq/IpDIF4/WQ7HIo90uCEOdH2iW7cjuu7YUDYnMy
Vlqy4gBhqZfPu8RvTAUI0i8qpUUrEoYhS7O97ZlHxlXYf+Q8f3l85d7fBFx0Lj0ol3NjD8G0a+jg
0qEiAwiMhteBY7AoadJV5+ZpbYhRqhrDLnRhPuopJAZli7hBVex8cLIoJn7yZj8S/XGuqiI7jJk+
rIRwfsdBUJDF/b04MX26Y7i2JJ9Il6+kewxw0PZry2QILDdmdO959N7sL5R+cKEO8fXcYwGLNGFR
zdpOKECJ7CHQNXp2yEhYS7yhpFuJQ4bJLfT3nnuUYZa1Urdpx6YqC2Uvk5UbM1ZlSuNx0c9k3mGY
R/LfWtrKy4b16f2ccK8onYhoCruK561WhaPln8bbC1TJqZNM+luaFPrzWJuw1nusWuQbBVeY+SgQ
I++L3wFqKiZUTmaeFWvxYh+Qa4wSEKqledGP8f+Ro4G3uD2RiVDOLLWiPdOyPOz1aRkZpdUU1Rcb
IDVpZnTLTakuEpiQ+lAIWLSwAp3AfNWawPcKr4j185lK/UHREZEqbejGJlLOEW48vzYh/LesMPwJ
hMvOfzRlHkuXnoKk2cyl3HP4lqMhknYIdsx4S+sXtOBRv84hXN5Khl1sm5rsilPksU8OyRVhZL5I
u01V5VHBvIw8ymctoomngUWvO4zIh8AkZ++a4VDjWhD8VOzI8KKrQs/SFFzjT91L4xi1lHnK2NhZ
AvIeg9KKmrWzHWdlWAgs0FyqzHvnEw+Hb6Oajww3vmEzqArxQdG3ne/pCXI3xpCQ617Vxlv0LiHD
Lf/m56ZREQN4PdYh+XO/a3HMEyHDd7GxIPLpCNd8C6zfXQI1kp96g6BAV/PVDtLBg/UEPObrZ+Ic
2thj+B20BpGX5re1ChErY9uBL+x9jNP8nW9kCkOnH193JhqhWdMicOQsfmR9bfSYvVuRpV8cirAf
SgO60BzFsIMZBthcu65SRpD8Wc9zXwl080wre6CDnpNmXeTAVAA+EcvnbQCno7wnrxu5npPIPlck
RY5J8k0BKBq5J5ALfNJNQfdPHHf53tm1q10naWSx2ocSMJ7xGGb9jwePhPVKPhsw8aEef0a+0ZNj
/woyuePqPwEqJJDkss89SCxpKKtWrGHhBbhhMBklqbrh2Wfm6fte1O5/DKOAuqqseQsePu3j5h6v
3E5iPKhsTJBwSCN9C1VLqFypqtDxJynv3jbNcnMrkakFYjq8mIvcFQAYUEW1hAsPFCdj/WEomDQJ
fyph+TSyzd2DiG0C27KIqQHgImDt18e9vQlXOqbSaSR2FasQgV9W6Pc9YfDR8beW0MfcbFGRaTqN
zA3Nv0MpOlZ9RycHpWrqM2ICLjepIoFNs776WSMuQFi5WNHZ+g3fsG5e+pQEQeq48q13pK4/qRT5
C0FWkeLNGw3sn3Urwm/O8R94c2FD7siJqyV/HjdZESj+fRqOjG6/T6quQKg8ZKmm1kO03CZVsWHi
QLxvFM45i//AeYhQI+mZulHHfHYutdwLY6qhk3A2L2LT4RNSJeZsJ9HJswvYwBuF9vWss3nb9ziE
uxRv7xqwNL9OL3D+dNSXa1k3n874qSkgRDkImS1fUKGkgyCAV4K5LzErR7HzYogcCCGAU561By0/
p/PiHVKfgwwiIrpGwXXSdeeRujlVVjmEbDbok7rHe2tYHQkyxEyYBsSO2miHb+aZTNTO96w49s/t
XlztLM/0eB6PNpcN1Jmpc4CLMmz/4cYdaVUAaNttQybaN4Mme3qr37pw4RkkIcegC1+Hay+s9pfO
URKmdy2yEXay5uG275xhfNrcP1iX26FOWWFWZUBtAJXrCuXUd0zJG2fa6W3pwci45292PNMjNa2v
PUzrEU6LxlIBybPDeLFUST51Avbyv224PFvi7w1Q6lYJt3McSoDusNLhcG859lnXcKxjU55/tJti
HFq2MARs+O43Xo1zFtjuPPKRu96PezMk+Ot7qfM/rNWf4LY73bDcoB1ZLg98Lr9qsyiHzfmhQOi7
QMpdn/1obn06dOouEXal2Ybw1SvLapsdOo2VEwN1AP9tQXPKTvpkF3OsThqA6EzmOY7i//RnjqQS
3rJLkhaOh7VmmQXZs9Lfx2rqb9jxFY3U4G7GvF3FoEFk3MOfPMKSuJEbYvlv7rHy+RoSp0vjeWP7
G52mq9pSW9enTwgR2J+2HALkvJ3V7VLKUsrYZR2SblGec08l6RKtn7pBgeXEL7S/VCxfzY6idGCK
o41atTetW4FUY2Vez4jBhy7EZkGnmwgoXWSwAZfUlTnGFjkefACnBoWLPWKZ2R+I29r5CFzMU/RL
EvTE3IXvA98BSpzXsx61YAESEProJnhUbV0vwvGZ3waNYNKxAh89D5Jqi4P0vaMA8S06fUKNFMmS
tjJeyk6Rvr+ZfqMxRdz0zl+9fEwiQuQcqz+zBQIt7J8grc4Mn+ugtQb6NEf67hniurEgtFG9KVXh
O0SMb13hVaRexNQl235Eq39CZGh5xx/tIF1FLotcosHhTL1JkPScBgduw2kYs38mOZkm9l0Gwq4x
EeifzxKzsj5YiUQe3RRYF+d4MklkimA/5drlB+ou+PbPipEJeQWykaWHQeMKblOCSLoXEm+jyQDY
yWtYI4tAcHnRM0TRvPKWrxglmo83JohFycCufWBELNojSPvh5Sf9WOzzWtRW6vYtOB71POtLLlhx
1mkAC46h5uEVlGvByyqi8vlGmSY1YyOZywewvc/z6EmEdiJLpjQ/sfMjxbLKXovBCnl82G5d2dVZ
9Kh8TCDMGzie7Kp+SGYndqvC9UeCyRuwN7QLuIIo0Y6jXha/YN62CqJa/jo3mgr6VEScqHZ9hZc+
cJ2Y1HxT3G/v9J//IsiyTrBtXgRaYzTxsrN+gLwY9SvEhOeNkI9m3Es9nmoz40Yv4cscIfELBAmd
O5v1DPjUAZmDvk5QH3csKypdxHRg7CVSu0jcqvZeAfxuh/uUwnrtD55Fb4x16uTso+LpF9aHp8BT
p2FsCyflv1+RN53XlM++pARV3wGCJq4xN3/UeZoXGxLBzyLrvuIxXMzUp9yCULD5tf47QzFNqtjG
+sDckoFCmtY8ze9vRx3s25Had9pUySOYOtxMCm6YXg749AWoZQrlUbuLazSyhIRfjz/1eFMQ+yPB
A9x50mNIS6NdRnYutE/GQuyT7p7I0H+TbN+OokzUAyu58dl5HVs3DINgLVV1EfOUQrT5hiyYxtbk
ynENtMTpZN+WcHFSdOk3fcEI5+o0vs8AUewApuzRNB+Ed7g2lga/OuLEOg+ZnEk83iIbRUnmjeXv
SJ/b9hBIT6Z2ksnJ+sKWbV7mEuw62RT8mgbVqkV2b6pnf5X4sQfyRl5LtNN8nzDq6VJU/osccwkG
wUSZvA18HDFnN/ygRwtCxwjq2R9Q3eIhnll82nsUnFnxuGFzFW9amDscLT3bUaBl2J59QhsVgrmQ
UwXiwEQt/2HH/kALI9KEWAnIW3ipN1aV4xKWq2Uv5zFIsSZ7o0OTiCWNw19LV4/n7Yk1G5IBKdli
QIV36q/XO1UFNjneBSo7SR0fBd8sZ1qSkwoYnOopu0kmFW2V7RG+sotlMVPHTZf3gE8ZcDTLKycH
8qYwWlqEXuHobN9OVVp3ciu2hppoPny6qPjvWYIclaLxuCxZqAUhWfd2ZKfBGHS1mXPpM1ElMJPG
f8RHHzxTXX1qymYd2g0mBM8twcQEhR0V8BBQfG9cmxyl7HGZA99aRhvGC237o7L2UTLoZylxjH2r
nTsEQPhLVDfy4vTHc2gJIheG1nWbZqbloBHWA0HYkBQEp6XZ4+V4wZKEI55C228nzIS2Hpk7grFo
umoSdKyhg4Gng3C85PTAFF7v6gwVhhHNm+EdDm8KP8xAYHFEbBxgcNzlNgsjGqNt0fWRPF5gAUPc
xNe5uhD1fATVLh1P/tPvC6qXryELyC7vsC48bEl+oxODX14xVxfpDcjFTTUcIoNVFVBqHi1FdrCJ
eqgx4/w6JQSBMRcjVhrT2Lt/61ZR2baYjHHI7e16GGkxzQGndQOUgkIlDW47X+LYtSJZmvS+h6XV
sbNG5rHa90s1irVdP/tMRllOLfJv9+1bixVsi1dPZDO/u6Ysb9zPjLh3/pXc0NRNbyiCeF+WAMLe
2/XS+QUXLaQrPF+ZgxRmBHmdl+XLs0kPc6p2U19aEqWZNml1e+Hn/uUQFbEpJSX0Zv9osoucLbQh
pmMK8DI9vrehg8CY4w3MbW0OGq5NVs5ZZ4kOygbANsX1wvO6CePQAelPWSAsResT9sCrJTfrglKr
kJJ1ZnyFBmDtft71i9R4AaePPvkMAiLgs/oGrhX2hAQ1ibHFNaUuR3QcRGXn/VcIHJXMhUZd4ymE
ZyPWgFbCncBoQBm8WIaZ+qwjzlN/wK0fvvSEpHIEZI6vmW0a9xiQrX3SNZOF2/7jF0P/XKDhoxkF
JOJDis7Sw1eli4gytKqf2i4hukjd+8xzVIcdvEiFPUddM+3I+XXuqmvJgOH11n7JwJGuLSbEjVef
rOcx0OshnaR+19g0umt2pGWUPFPQa64wM/b1azS/Zn3gW+hRvqRD3qteijPLekuAHrAyJs8/Hbhe
hl0Y5OZQE4bmd8uewzA8RZdSOY6FdZaCBdBkJFsklcinedGJMjp84iwBCG37iG3UnHHQU+4ABZIm
8Jkn7fCn9THEKsmFZfstQgMWtRejBkzpbFIK8frb7c53Ms3aaw+/xn6ZHhFxMOuW8nd85ObhAvEb
z6AX9lnrpjMdYlQjad9QgevXy68sue3w/ddcHOQ7Wao/7d13N0tOUByWZxRH7k0cnJuGrE95oN+b
g/Cv2PAQAf4DqWhFUFz/FSwN0B7ShbltAz6eRLmP4fRwVegprh3MknC4ZRnv9OsfVzPuRC5xO3vN
SSb8oJhUFOUNxR8/o6ZRWLhMFpUDHLsvw/2kZ3nhz6826XOjA7wnHWwTctSFzrnjFvtacfz368tX
gyydnjP5BMOATg8bUAJ3Al1LoOlNRUCOyDLjrG9Yy8lN8oczQyF5WkaFxmiELdZOhznrdZM9e/n4
j38QJlbpQfqhVQamjeGJ+VsPrUZtcmnC9Md0XIt/cs/Lh5nkxaeRF1kHsHQPwLnZgXa7PBeq/dhZ
giCnsueR2zvTzKnK6ixQEJ3gl3jbWQsR/eFy4ufxY0NZzmkUgpa8iej02FnbdfjSC+pzvI7sf4QF
bgoP/XKZ9vwyY+U/BfmQjJ3nzz0YdjiCLUo4LWWbK9Xm35afPb1NKo0u32+2gugQMbNW4JwQpzW9
G73u29dca/G639ct0dFjC0cKkg2b5bFz1MC1T6j77Zq/MnxETsaXpsnet5nHxNI8cqNG0/32DNO0
+563AO4GycJZPnXAkvD9YXcuL2H3Zc5FneVhZ/M4r6Q0xuULaZHbRS4gdEwK1phJ77pllWcYu1G+
EJAG8Qn+zO5AhxXhDY+/Vlm7nlYaZUomYJqQ/SvKI97xTsayh2mIey2eM09tqclT2YFX5LvVGda8
v8DfG6LWHJWjbRaE4ZB8w2UvRsdheFQvWvGd+Uy3n4kHv+7Ix8AWv4N7u5fjRSkWOA16EEDZE6oS
e88XEquZDKU6oskVmAfMpohQVEWKmq2D8KpTUwE73VMtBz8HuvHin1ogf2bHFANhhgmif2B44NTz
tLgYwa3RQALj6+73DlnJ7qLDQNpFnKpsfm/+VAmSGOKKR+MK0hpskEofJFUleFNOX0cuaHG/AKWo
C6xMtMElmAIjOoB/5UyKAlzk4a/HqKmUqB6f6gy550/5IiT+GLt//skMVb+oNmbDvQCzXMcN6tvL
sywocmtYw16/DU1COMAnhjxohnKfnlnOZA+uXEmNt2u0eyhhOx2IYOOmjOaiQdbodOEbxvxsu15k
7WaBugTsng6Tx2Jk3fgjbzAcp3mm6ovJYgpkt618jDbXCa3qmSY+fwQU4145/VsbrPRhA/jQ130q
bba+XDed9gHMpRdlYg3OEPcVUiXRZQHYQv3H4lMUktlccHtgl/js3GcupXtvQGV7D3N1QHvy/BNW
YLBMQA7vLlPKFmOQd2HMjShHtqDtkwuK7+mrqzidJcnvEte0oVZ+O3spBDxJjhjOspjFdfxTKa0/
pQj0bHFuNUpA5WdYX3ct/MkcEo6T4tgp3jHjNyUff8JfJLT4UoKC2JhiLsuP6chaYmiyC3TC4VQM
S7nvdlo1fJ5ecmE1wG+uzfNxBOy5PQvHOGMnH1sTnHrZWZBznlIUIrgHr1TiPqMduSnsoM4a6k2W
+f+NN5QAASgUY7F0Jbhbpilz5rtvNEvPBUckyAycRWiDQIrDccFo9FaNZ3aUP/M2275OTl5ruQi6
ybCobhEwWmDC1+SG8pAnLNdV8NjpTWUgzm8SdEN3SbdSh1TC81NMjsEqxWZsC9x/N7HjuzIZrWl5
QDeKeJpZ8/ymmOIm2y4U5OFcohVtEwAR+jv3Xcgxzajef8jFXwxE23mvDfDu/T6t8oyfvYjvuE/Y
6ySk+fMHf/txMhc28u/xjlEQyksiOu8/fVQuM82vdAg9eudoNrPezinFQ8rzL/K5mCOS6yYieLt/
3owOu7EoIN65IwvXJtZdkz1Fcf6jyCAzXXuJIYWLM0E7u9dytwRcEWcFRCNJGhpr1w1c+heYWTwH
ZWFfkcJmE7rNn6gM4s+kSuQts7qb/gP5x/qO5vtVEiHcSq+im1Rb4PlD8RPlHc7kvTvheaf+M77C
2X+gMt3RF5ZU18hMEZ8QVipLCl5GNgJ5XHrGcch564+WJXCkKj9xnKESKYOC4Y2R3Dtdt4/v4gSp
olhAY1c3lKEh+6KiKronm3yENot98RXWr8YLTARUzXcn2KmWQf9BaeMu8RN/xEa79u3Xdl6fQZFA
9ylnAxBnaNIuwiYnCM9HAjFPefz0Ax5C3ATs8jC0pLFDzfQEmchPFg4qJWndhCbv+JbXjR8IJ62n
ZIR7zAPViGJXvGGw1hUQmS4YoVkOAuZQfKx5UtI1xFhLJBgvLCFybPOporj26lN2EwGt9ztRl4xC
vHpAB044FwcLmHDppy4KRBEaiCaZiBs8TRSv+nkV547lqaVrQgIZsk8ZgFc7piXtn23RgTJV3f8H
2N1VDvoAINfD/JrODtKFYpoSe0SbKAipPMJTRHU7IV9TK6302lbP2wK3FgDelS7qDnA8li2jOhCS
CptNfhXpNDlaeKGszdCCTpydIETNwFOVnecUuB3q7SuZFh5YJyoCaeDuCTbNX5U0W9feTOpipHo9
aYFlhwW9lqRGO0vJmcj89xGVhj90gfp39FNpZL34htEvXxxCpJE+Zli74g+xHU1TsdkGOS7pMJzu
HmFDLdRHIpwlOFkp2Z3KUz5yPvRHmYOJ6mRyoV0BOA7kK3MurC0Y3fdnNlN5hnoSlA1S9iPZ1Uwn
/X4iysm4eMQdWsCVquKi4nISIU7DGDhzTd2x7dpLUKTqWYPI041fOwk4XJXdgwC1laVoPekPytyz
bCGZlRv/OwDQ2H4kuPQPrEamwcW5a1L6oauh0c8ty4v6W7ANKc5NQuJ5pqQqnJ4c7nrZfc0muZSD
lKZwagjajEPBA3AhO1b0KMIVj8JsMofp4qb7nt7e5TMp+O0wnRIOWzzZKcRnoBffaSQYyE2S+gw4
izL7Eb4pNWKNV9g7qStfy1ypZthPJJMswh6oSV+2DNgrXX9aOu65Vxih6ygjRuk8yhh1oSLcSNwI
7Qguidv0fiEemN5hjzdSF6eXVOovemG9CnsNCRDx5LmtsyIfn6Xh6k9yOo7UAvyVv31imuOmr8JZ
qXk9Rwtsu4fc01/XvedZWvbBiqmduDE76mlsQ+A6XjtqYjjNPd2mndfvxs093d/Zwu5Z1iLTiHnB
XJd3HcHbIocG3Ayjq7yebNZ9vEvgTRmb0B+0Ph/RsfmJ5iZmGGGdytSfdaV8ppFsU8DdDdOeB0bw
3udeOTh937xahgQGGUp+pIfrhuDMvMcHa3kI/WBogX8H3jDoUoMzb7fMxYeZQBgUREj+ZUqzTujw
FGnsfK95bIEui5pyR1Jbomq94/8wxw4YXcCNwy041Do27Dpi7wL/W5lt3eZzJwjyexJLhXzevqLH
6GRFhMi1Zyd7RY/1nlJWX8XXyRmpl5R6hdlG8xETe55ButvFJE+BJjsE6X9ilVdErY45wd2ZiwzY
+JrRLth+qjbDX8+WYGfLObjniaPYF7zt8T5Z5f3auUJhL516Lpw8/ug9y361HzWMDYqMb2kvMiRT
+a5mIIJiT562SEWaa4UH++SpSqPntTIejg6K0Hc5mRvsKsq9oIOqpG1Tai3LdMN5o/4WKHsWr2Ca
gW7/2kNdP6UUHFBzFxiOk9z6Bu3rfKZL0bphHATU7EFhIrQPWaa5lLMBVfNtUzymIKSG+syz/hO3
GMrvuJSLUbmEZnTH5obASxH9NUHPISHFJfwmQ/0SAzXPXPNAqfFl5np6s4xXBq2lhOXd6FBAEpWg
JzFYWoXFr/KRCQuLiwt64MUzIVY5bRqRx2CpLs3l3TnRKrZAo/MeF6O6O5/wpgDz3zxqTJo/hODH
qxNDfoFMdtd8zD/e/42/gXvpQ4MIaSuHXH8siQNcd1c85gmGCTF7Ds2QL50zIU4o0nVirZYGhucO
aReguH85CvshpHtnvMMh/e36ufO7ZPSmcAjqpyKgorsCRwG/WZmQJ5JIZVyDbPRiLLnhjWllywF+
yQgAJFI85Z5FSBceJrigOnKegW23ybylXeJz2Zr/6Rg3Xs3a5uMquXYBtL7DF964yGdv+gSk9LXW
U1g/tMVz464IgrAJ6PZiSaE0AkZcOHqg82UWlO4eZs4Vl6LaGYnHEHNZyUIO3NQXgeX4qKQyiVqw
RPaFpgS/LXZ1WwKunITNOc7VQW0vz5SgSONi7tTV4BG3g4/YtoS2cES8qTqGtgijzuVLYqnN6o1r
DEVK02jO6I5JjzklRe3jNXuNwDwDfnoZ05GtdlM1EAenbAb5/Eh6ryAqpCPyj/xKT3nOSbB5were
xeBpIPWsMxGqGwWPRLZlTpvsTzaU6eyQYEMZIqdcignasFJj/F9Q8+FhjATyFIrYQICRd2/noKUU
4xof044TevIdCSYDtXOwWWAey+u6ZlXvKEFOOmPAtvKgh4eNSuSMullC1zdz35ACLwk3D8jQhTNV
7n3I99v0jySw8wuvVhPNh+styde5HCG2TmxOUZjYWS7PjNUwlOOy41HgQu2Tj1a3hYJs36pzeILP
oSYEFHj390+hvK0ScJC72Ns1Bv2XR73VcIOCzbJSxzLP1HeHNrKf8RDJHZWWmPCamXlIiPmjqAe1
k3VT3IxfsYTakhlNxsfc64+qVHkfv7kS9OnATX4hLzrU38XqbcXxZj7+r28bb6c3exaHmFtcJtql
zJod/1rC8NWXhoMGMET1RrdSED7HvtI5FePfXqZQpmB4z/8WogSxpOwzZfecNxzv9s5Aa/RnD6sO
8pmtuXJ+x4CWEofgWFF3DT17ouvSbmiizaloCLPlENxisAGlA6cf367FgAJuhA/gz5oxBMiCXcKZ
DuHw12ITXjcgDNCF4byb4K6guG+NVWjmknvfaEO5bBfjWRlvVT8RuB2YzWKW63GqvXqUa1Fzkmke
hM3qAxlIeMQILTmogCVhPLDUmWN6K8SO/tRcD2uqsL2qE3AzEBJK/fbX65c1vMYB2om+t1zQUAzO
Kaj6LIyxYuAq51D4egdb7+dcMdXATmzOYNecDEaasN1z5QqdQHb/oYhVpB13pu1lT2ysinxCKJCV
N2gjCpDCh89MLAoxuMVqmGyyrICdTCBnQPPkpcVgRs8jzjePUDkRgV2IMstPXLPkXN6A5M1uHJY/
jhOBdmzYgQfpj5LDqe7sPH3ET8zoHvxXz6912eSMlLYJO/VP3CuIxtQZKK9j/3wtTELArKVCFPGS
fRHStEO9ROdJo96HIwRzl+BfnPW3P/AtDIjxnuLOV05CyCXsQQkvurS362T1RD89CRCNiZcgp9uv
fG/47anRsaozoxxE+dKpTKL+pYBQl0zOZdBW64lTvc3BFZ1YOApt0ZpqLa1pWng24HYZ8APzcRkk
xqIFpPANXZvRAu4VgkLmIb6lYshezpQI+8wNSTABnrlyLla3ZN0DRGZ19CJf3PhzDPVbdhEnUPa0
U11IPihUugT25Fd9Qa2A6xEqD8/+df2sNvelt4ilSLiOd0Z083WX0wfEvIX5GxOF8i2uUFFEQQ3B
mhP0soFCNOSB3M7vVfpZPSaDtHI1GCLGTTZWLQLsJ+XC1eTW3fCEQecmMzrLTow9qvBGy3192Aip
TtjAdTQG3dzMFmMYijBHIt5SCOPnoBoBe+M1dNhKoYT6iupQ085YFh8qexCVipvXyMucoMgvo0Da
/ogVBND+cwqqp/fC5N51/VWKo2tFGqvz7xdx8CdpzgaUN9jMyCuu/lNJNERkL/COb71/PbL+Zg7O
U9FnnGTNptCplQAT9+epGUTnfpALIUoAqNUNw7aWzm+lZDfs2lZW3VD/JxLEN88E2cUX7Tkbq28I
BRQMLhskLQ08SqnR3RfdHUul9kcMzR2Brc4ZWq+/EG/sZrVvKasy6KfpMsPpC89ENWUjElw3/okA
Q6dHjhCpyaD7fsr84bMBHqVhRuKWp5/Beq5GGCjmAFZX3unkOg+tn5PvOnj9Kx0BxZyJUP0T5g99
PwxcwQEUmHI1EWxJyxsRFvIWXzxIyYqtIJsBATSCWeM5M2Ad2vUz6yn/uqc0lsF+XACzk3cMQlhQ
+AElMNDO1BuF5BElnddOzsmdABn5sPPXPKgtdgFr0pCRDB/1cHBOiZawA7TzoLzcElAvQDhBe4bo
iI4pgvJrSuku0fCzLAxwFy1QA+FO+yrP71wpQ7FqAUTc6UtKCBuEaQqKsp/Iyb3OIDrVg4sGQpm5
0aBtoKZ3nxCl4G2BLLd5fjy+YkdfxDXDzbMuw4c46zb8qfJdV8WOeCOexogwr4VC+nVu39SqQjK5
etHTdPe511mnX1Q0XCGrEDCEa2vXOynsUmev+NgRFqPsavxdCrFgKdm5nOzfjbzHHFXYaoQ2o1Or
DAemAdxAz1pdKfVLPL+/QzHEc+E7E7KwoPBq58UsjssiaqwxquR11MTlAiJUR9Xr2Vl1uCifyeHQ
3b3htJksuZI7wPnJieFUnGUaZBr9vSd+CpLsM2bz0hwuT7OfU50FHJojtwv/2+2jRV7pFaf0TTFI
kyW5igAOYaUustYiccmlbX5cn0U+cfa1AKAw7l5odm80nLgDm1+cBvxAAhrjy+oL3XqHzkeHX+La
kaJF3NfRyo4QVAKcgCgwH7O6WOMipUUH9LfJyUyhSq1lTh1rEeup6uAOrmJCTkCypZiapR4qr69H
/OzzOfRVgTiYvXeu/PICX7zFptr28f1oTc3ATk9NNql1rvq23Cjm0cPIZziI69mYIv2WEdM8YWC5
0ubnRWWCbX4Cz50yY5Tnr7GKR6TbjMPmM6g+XV853GqztbUgl+wLtywsdHbKozpHmTT+swwkxJTf
Z6MPmKLhEM61vIvu0vOoL8qpUezJOvo/BEK/oztIXyXlPGrEfYwsIqy4IWSnGW636DHPvIo9Y6Ga
/sZQxcd2az6Qsih2dSORuOu6yxc51KmNujfeV6lDXNIIJ70Zk5ydjj0Bn+62cid+SiYHuyRfofup
cDU0EJmRKRKvOVHhZzxgPTpkzPiirW3OSJrGd7gZFAZz+r8M9ocFVmJ874F82fcIN++8NxXPgNfv
EwuPj8gjx/qvJZKJCenRTJY0jM5lLx+CaOOXM3Ww46R86VhI7AMlYak0hJ7JKaNAYSnIdOqFeiEr
JDfw5pCrMo2BHLDNQu0PQ+ho4v9ZoMJwTS93MP1aI30nBUIkz/VTryOTea7CZFB/a92WV9n9d1ox
TTvETgFgCbLFlICFLKG9rywAPGa3dyoSeKo/bFreiVFfTCJh2RZQCokHE39NbPk4sBlOi2LkJrmd
D6yo41IzN1cx3IHS29QYS8BYhCpjOaxh+yqWDB8TihI6KeMP7CoSRWTikn98Kz0r8b8N9y47sH/V
x9RiJNbr11Wto/R7MIt/oYPPqwA5IqmLMotsdp2mU8vcDyZhC1LnTlRvbAASmIs1DUeTHtcdyIP7
/GVuuTUZRQ4YnUy7RwovPVQhhZk673BGzB4VFaERkvYABkRTpEtjZPTvwhuVVoEr452/wUyv3GOc
BXcUET0VAf40fcK9nCHyyVPo/p+UgRmzOvHz+B/3FZhkaGC07eiLCm1u/Odl6mE998wdkar/aMKH
9MsxEndPdZG62un9HYjLAoLbPBJjrCbGTJ4GwfjOsbFndMEA+iyfhgqq2mE/tBP1P3QwaWm1l+Vl
Ry8efxIq74WETAVPPTYT3IH2AjL7NQ6ouFLxJHgS0sWzTmLqC8OtJebQ/z2NoSYZJEGA0sRiM9G1
RmyS3FOxYTx/y3Hxm1zvkAXhD00gex1VJhvEt0ZwFMVxHTtiPEanSE3cqivyTzaxLx6zqgI+c9Pp
XdyymiGc1uAE7PK4amturm5mxFaTzoFJ+0oqycIqI4Kst2xGle4OAl36kV4WN3lHeD/zOI/6Z8Fr
PIEkcFTis7aA8HKlqYTXPeBbLMhcpv5G+hd5Xg7RAooVSTqR6XeyWoeuIZ4qcC2I+4fTHvIJzbFP
3PGwL2tXSM0YajU+U55Ftw0H3dO/jw0LeEbzEKYv68mmpQ1VblHrw3Ta74uak89XJyIwBAa1LZCF
T1kfEnLMMwnZGMIvKbzXNGikJt+0EK47NtZFWX9wRo8bkG3eZa4h7Pjnwqag7SeY7zRMxycQC2aB
PeBVX48TP90T4w0juY3tuWmC5nnunkBilJ+VAUkwQH4oXV+ng6XTUrPagRZLMCpkAGWh85dO5AJw
sR+Q76NYp8vgC8JLpZhVRQh2UBOo23n3HLE2w7yonvaL5G2LgkDEoUJ6tDl7E6Pom3ZtelQFpgDk
pWhxLSwz814yURBM41Fh9bCc8cOjzqUgDreGgJZVx9BhMI/+OfZpNF3kge7ngo4hVYikqwiB/EBq
2kp0sQ3sXBO+L30CiVjva5inP2aWjjYNco2qzljZMQLh3IWGQJGn+QlgVrZQgJ9rW5br9hzxQVc8
psaPxAsqdJ5wKfjWfoR+zWteKDAjbOlUouw7AyBlrL+0tykSuyUvQ/cmLPQ0qAnG+bPSVuWsrajq
5P72FEX5x+pqFqtSh9J4zYD0SJw4gwCEiWjsLo0K4rxvWnGtwd7wVfq1gM0FSf45AenvNChBi+/E
0+4f7kpm6XLULOIdKet7FhLXskTx0L+VuhNr9Gg6LUXWIdzpF3BQSYK+AuouxlVepVOwGNGTcY08
rWefbefKNdGfyp9o+gNerqH4xsl7U7P0qieU5VfC5WImmmB+vkdXjX/GN3Yw9qMquD/OMUY2jTXK
SjB2Y5+3C6qPbZEXysO1C/MfoeFCZMe38yCv3WFnlrwDs9hEH/EzySRpzQHIXN0jPMA3alaEgyxY
HnSLoY+8iVbgEEYj8I6at76mcyYbCehSAu3nHJWuZe8d7lQtDXQY9eyYI8uzoohs3DIMYznWc4wZ
5Ga1W/ZzAthgruusv3c4Ub15xWGhnxHfz2bH2lYVOsGaD9q3uQxGRnoRdT6H4a1PQFud8yX/ImRz
WLHyGRyuRKkYif6/nAxOCxE/HTTMIubP308zNGLkJIELxicfz6fDfwdxsuad8UgUn5kW13jOgzKh
d8racFP9XL5KUKAQsSQed55gud81yNiJPdWyyhlCdbBtxDp1b/cKLHzIfQev7SwlqNMTYvNqAE7w
nAtQcNMK00l4Fw50cQNyW2UMcUWZlqrLHYzvGUWdNDq66vnhGm4SWqaKqXttqs+TIYch2AhUTgQL
rjXzt7AHnSQkBiDdpia7oV1HbkU95lpaPEWTOyujBsnV2YxZc6gk8cM3THOtVbAb/8oAN/TGmcfT
4bH0LGBszna/9FRHWxN/wTDDsF8SL3MC5cy6yMGmaOkWnlcrrG4Oq5Xjn3HPOXGNtQ817N2Os9Ei
34Zdd+irQ+Q6xx+0dYF8+1uCIATfi7LRzMoLGkfMsveut919tHBx3U3nodXNBOZxytVH2h61maNZ
9t4ovITnIseEuOxig/m2A84Y4ZgxEMq1DMQaUDc88PegkhtPVeB1X1Wb/DIhAJmIXRH9WdlXvCqY
NdtfjGp2xKWjb5e+2tUxJulPEoZ0IoKUBzp1YbZP+5csAyfBrKJ3jeHC9NYq/KsoOsAKFdBRVUo7
Uq1WCN2w/Dzpntnyt5xC0sycpOelzCyfT0wakQ/E7TRvHx4uQc++2cuje7+triPMO0LrxKs9Jyti
fSEq1xIY8L4oHfqv4xIQqTak0SnhS4vrukE6/IpC7V0ttJU6mPwRDNJw5ok2NebZojDGtUZj6i4b
Xc3xMnDNIh4Dl8G4JKuHyf5CpCItwG1kirWg78WKeAKOnRINq9aCwLTYmGMOOELzqnmvZPSfJIJL
BuT02+Kj/IoS9f6L/+V92Eu19YUACdcLA9l0JeSa0Slmj71lWnqtWHtrQxW8je1C++yYkS4PBtBb
qQlOrPtYNxiCgYpmBUdT4Zsi9mcVhZUHX2r2JgjVEvJOwVze0sUsjHKGmiOpmymGmzrTugdw+z+F
qlZHgjRTIx5wuMO7VLbK0khUvBbrqvCNXeAYyK0j7wc4VcI18Y7pNFTB4Ra6M8uHpIQ6oHxQqdA5
PNGH78LXsHMlgXYwJ0quNZIt2XPSFndR3tfgQsT7o/ivYGXdRjtI6woberkR+cXyINmRQwZdWPNT
er7yydT1wf7Pe1jDY1Wvld6jeAnfFoh+6WGTcp8sAMtBQpfkL80zck0GEP+4/HScfDz5VnVKVsu4
702wUQL5nf8Dkex18h5A9nDcY5MbhqdBAO+e+KsKY7i5fWp3FutdNnDxn+3WTYv+BL9P93Nvo+M2
KrfQH0quTKviwPdgvnQaaF8zneOWWz6J6AjEGoFONsbtHBc3eeb4V1vakLlwRKAqoNDaizGjcrCH
5GrXrxAcbyxDoPDsAUJQNrDbznRi1Tg4wqVDUwZQsmE+Vv4Suy2vAm0MIUpqkf4E/8QfW8LHKNNq
kNcHdm2vsAkPMOX0EOQ/sN7cQ2EjDak1SzFWxcoe7Ur1umtRYY0oOsPSfXzdwHTcd68bLQw73SrM
twLIZC2NGfdueS937V5QzC6y8eEX5k6AUZqLYp81v9ld3Gd14hjsIqUage1LMV+VEz5ACdsMYSW+
9grCEbd/jeLLsfx/aKwDY2G8j3yiujz2oRpaxfxV70ZBfvu9BrC8EV4T3PqKAlFEMD+HnVHNGNbs
0LocuyIzzeEzKZf5BE1DBs1vuykupFTNmxXWmJTnmNJPKGg2Pj0CpKPWtbIR5yDSgegzlFCtQLIH
8hq5VxwO5hpGyP50yPtzFh4pv8cvw5Br99ky5ovi9Hx7FpBy9ETPEnzepz/86gTaBxUb9PdhoQFd
huha6cLaSiOK56dWlTKo7h1KAXtHnLLW+eKKfO5PQ7kOvJvfYew/NtnRomKn0okJWIOLbFYqnLMt
V/NCu+Jxis0sld06Ij5YrLhL3HkQnMthP9Rub+1EeFRIlNnDX7LPw8bPTSKxLLim92H+7rezNjbU
S0SGgZSn31SqXmGPeeGJ9LTGlHQf2lPwHGUDKlIiOj5N8Ke+58SE/9R7exeOtFHxDyM6iKay32ga
d5CaaP6RJw+QL2we87Vi97mdjjMrzB7m6bW7ypXNFQEbkN2QmooF0oXOa3ExvwMxcxFGqAgMTLve
UDaVjDRo/s0Ub1gJJm9ebdKis+NzBZZ5fCltglv/Ey0s/2QR2q8rq4S1ygR8LjjvKoukvfScx62L
4ApMVli8dAK99poY6I8ufOuKGae63tX/VrQmwzAOOGtDcIw39f1Zm9lyZpRbnItNmIE8letx7zNI
BRpkiv4fZUvBSihFe0qLhQcvQWsIXR6n2QbwdDnSMdnsFiH7aUROEmYc5kj1BkcqcP3wBbevOxvz
ODM9rXZxRIiWLVVN7MFu7MejWaLQScPGcfc7Ybp0yxI1lzi9izJtRY8oVq0XJLCXnt9dYKg4E/TX
YqiDfNXOKUGNt0rExFbJyHiXXz+HlU61PlNRHmXaMY+s0wEtOwr4DLssKGXfLnpBYdm0ePMh4YS+
09J8qi3I6fVOHZaMgx/EQv/uI6sWtxtG8UgVnADf619zl5tfCJqITDFD8i6rdjDW5JJHu0i4ifY1
j4xMkdTMg6kKch/prW8+Xon2zbrnod/XXGn8pbFytfHRsPWj/ppFJfxDD8SQJTDohkZItpW+/fgz
Zt03pxj4JpBT3F+qMyXyU7qpnBXOL3bwnBw8ez5WzC3dBuWFTe1BkgtFm45nSWdM/m+FmrckOQEw
Bpo4CFt8orv4r2Bd6tdUnsKCARVXO1mucrfTa3RGlykh56Y8ADX8aIk37zAXhGfAwe+SA+qBiLIr
akpZWocGlJKV8Ol/beWOwF31jflZqzwZwqYYaZxdEAQuV3GDdTejNL7Jnc+ZZFom7Eg76L2yAGt5
YyazC/LWOOuke4MHL0hmniiEaYoOvdnJAAfPGJbB8PJ35QIIqTvT/4OOA5MsRffEKnPGskodh77v
YGjScHCcf3h7Vf7ECkZrtwjNqUSzX6TGvnK0XGsvqxVeaj8m6uMU2rLV55wefxP14dvMLapsSJ3A
+9P6IoKfk1OGr5/mYyJtH7DhmNMhKJLRkiVvpX3XaYOq62xG4vQoocbqByv9cPy02oPah8qD3Tug
M5/uDbg6vhp7lPxGha4W4TEx8IPs/4cfcsOT4USLRDzUohbGWrajPzq4ClBZ9jzhuULAu8rXzk63
iSAmrlCvsAvU1RTL0vvNwEJU4Gz7JXodxMLrzT0gZRDjCOrG+f2xOuiKGxAcWjrzJAIjrEh6CJDj
gz1vR/D575STvpXKw1r83gh4smKWsPDGdoh1Kys2VGse9a0bsNslVpKMVDKQXFpE7vcDSFg5+8Fn
t9wEjO4tyHZx0C34aQL36lwHQZRtp1VFdj1p5IXMYmK6DTk/40N5ZjeF+jIMsw48cHrnXwrLcVPI
JAxdCQstx6tCLDTnPWugkxys/oxtT+qEqdQK7JfAV0NG8eBKu+I8JRB9hIra1AecZxHNPHoxXv33
D2piRInUug8USoP0RBsJ0Z4Gjv3fRRgnThGuNmzYZn4gJBoIzRBnexDzPPn7dFWA+11t8sEAZceJ
FaMVTC8WjD+tJO+xFbdNTbvp3ULfPNEAwRaZHbEsWo7X6EzlJccGUQ24yeB1QOKwlFyR8ve10GKF
z8nkrFN9y0whKFlqNKuXlSV5W6EuHhz6igRS5sBfeorG4Ojon0Rc50Y1Py4l6OMyxVS4XrGiwHuz
I0rOH+cHyuNACkzZOU4mbQdilRUsEdFP4DdAlWBjNeLNu35t/OVXWQoBFO4XPFWsWdVl27g+/hqZ
U0BSsSGxFvesRhE82IEI16PPAsmTUhajKAg3mO9sRTPUMTBVREGtQnjA7QmHkDMCSmiGQKsE61D6
5nSDHgzLnoT9WpnBgPkjs631AiGR1duQbj+tshPgC2HL7S3+CxRdQt9QlB/FIF91CS7lp2ur/F5T
2psflxf5leAZfC11p2q5q9O4tJl5oUFQXoFXVNaf+lBBz2fRg3t2UQpOLAjFEIX2uf9cr6Qu9998
tc2uDuXdvSYYeAJ/v66NZixtS6O0yaCBAn67eYqtQY3Zh+PwNkL7Cog5WVwulzeTq6iw2zaTRdnu
lWblcBmn53eU+LQmvuA40oGh5ACQvHNiIJ6kL3sDNMX0u63PxWrombNWEvaMm6q2lCJlaWUCvo3J
T6QPDRmQro2uz6SID5VyhX+frEG0YXuszs1mPLfKMkCRoYa4PgDHekWq+lTu27Mz3gfQi+VJhzS2
qdZxNXxIIz/HQ7soPmL0Hvr5fGFEsXSbj0jvNYlN5KPqKuC6FTKLg8RtCpz/hpLsJAUrW4mobfPz
6GvMM/s2tDjttYRYHOAlUD2DGssr8OUnwSPZKo+BUf1HUBys9UWX55MaQKWow+n/T3N/2fmAZslX
ZnQh38oyft65zn7Bvkx1DN5fOJ9mKaxAS/55mvhWHNXRkgFV/1eKF0u1hFlcNCR+Gp/BLkbmY9Zk
9gJMNBsZfS5OVs9NmKQ1WqjbxOHkioj7/tC6aauTGz38j1FqCBRnfPJXb4rEq7LMmm0ARaz0hD32
otE2svfbNYWzm+kV2Ui+iNPwmH7uHY4jaaEo4UKkVeOgjg/B9xeyfMu1JJ2BlIm5N3D9Lg26Z3Xk
I9Dh2VLgJgJO+Evf0Y7jrmrv+v4NAsjUhLfBpM90TGtihL53NOOs0Z6ga57E9UbmkJh1nf+anMoz
Q0UPGtxwm1u0eB3O0jJ9KStRUvE7f2qrJItd2UmaCe9cyVdjFTqAs+u7oPD/7EZSu7Yb2eDgwzoS
d9VaxWPy6xfDMGz4Idc+lsmjLN6yc6qzHapEwFfypSxJ30EE4xx9frec58dhY9FAzt0uwATqUEg2
yrQ8zMKoxe7OzgR6yw75zQIEzcJCnpIeWBroqfMQF9HbeuI3XxF7T+R1olCQRh7uTb/hgu2zj9lD
l4PadzgoXxjxVQNcraK8+r+5NqxWsntaBatKgguJiNPN1ugH2M6JKlIuZ35DsnmC/syOfIsQ4hz1
2hi1HF26bawQJZDPs0UxA++Nw2ve4heyFstiLP51HNyEOdATJvKH2XGBDnzkm9B/nquJ9p8RNyHr
++qMdnL2qBzogsXxwkCpBXxEsPegSVwge6QuF50GnDN+YrYxeRE5/v/S5SkNZK/2skhB1y0p2OmI
DSv8fKq0NxKzcemGTKgZO3i0GOXe4zxuVgBTKqjLKzHOuKBGuBDBxaWUgmuzPBd4pkn6LIQkYzPm
RHmXRfgOrKb7ZyQAJy5M3d5cY1CCTbki1EI4iyZcujuTeN7Eo30dhrfYV0WkQglnYwGMdUPGt3aG
0U4AdNujYvJzDP7/zWAQOXAo/dX4ZFGLBlCUXa+mri2EI1Bp2L6ECXOVWiJjVjP371xRXq4ziDPs
UPKiQ5ycEYfrJ02Qi4tO6lc0LkAPD2WpyffZW3v0g3PRXzzKBvsD8vSB1GBtaN9oGS46Zv44Wjzw
1hgRpdf7wUlGML2+li6zjPfOj6EYSkctXc2+fc71sp7FlwjzLfYf73dojz+s3Q0wTMJ8l5j5o9mF
luRe/9m9Dc4SK6JLczC5ct5+QxylWQD1JfDtdgXgQAuTXlTdf3luuZAPV9FHf3/JpmmDvw9FtBlk
j8g3xvaWxKQRYW1QCPKwlcp9xrlhO/A10gxEayBEZERp4E1x1Oxu0S0Bjidwm7MeaJNzGGWg4Rsv
oduHbltj79Ojh8FhrE4tVG/ilImX4yntYlLx5uF3Hp4BpuXs9R1FvkRXYpsXg+GIt4h+pczR+ioi
M5tR3Ad4ayAbygFr73/LnvJlJ5RPzsgq6Ss+dxOwsvDGpe1r7J3ih2veW6EMR/69Nvp8j6b40u55
/Bm+yOaMFFcVQMWpZgsmzQ0tgho4c5F6UPE0u2sI0yPM/Q6u74b/1vK14FEzbuCaQHXMFIId3dub
oyepOwG/nxuER4gQqYPaQtjfgg0EumiMXF680f2b9/DaQrvoK3e+SceQqjGpjzQRfEi6HYokTs72
/3il2jMFFft+HxSgljT67/DBPbaCJ/iMHqH9mjqApU9wJhNgQ7VWpaprSTkwySgo8RZtrIGYhZz9
Xw0n/M6r0oHK8rohHiOm+U6fVJ5Rnev37N+fQWG6tUWGeNx7z4vMP0lNuBwnikjpnhkU+Z7wMGGQ
+s8GV8tNFHH7J9jadDOovGTH6VN5f0sOfGwxMuElWUU9Bf5kGVd80gUR+kJs8pfXSGuKaq6na8N+
FRrwDEGjas55NIp7oMFhyuqztJPipFfN9DSfpY8iY2FI6uY8fg7S+sCCZkOISbGsvO4hRjLM7zLs
tgQA8+oDW4ZGtGFWeYILIki1YMF1A9rc88svPhltdLYZR+pRi3mwPWVfcQxkC/tH/TvXHUpldb8W
Szr1DPEEEcnRJDVXuvTLImpZulLk+oJO1CyiwcHe66oIsVUO4+wmMZ79FleBgfDRKq0+erXcGc1l
u4uymU3Zf1qFpsW6pW0TG0trfpoi61fT/cC8W6pHOIx5thkC/cTDMWyaKy3YIEc9ueCa1F+W8QNQ
LWpOW/iK9SlPGzc8qYvdz5vl+WxhvHFfoKO7mO/8C9PcB8lroLVwhe3Vy1sym5PYqDwb88jxzNGn
epzbdVDmqjwlSfgV3DRIi6JvULy0mfDDgoBypBkYNTkGUb9CwrdXCGoshBJOSZynr4aZd77dlVs2
oKETtERvY58kc89agsknTx/kM4wkr+jFWvTLXDqa7oaHpdirnr6PG++MqYVxB4nnSbTo2xrr6a9p
lQ8Yk7Xu6SeOCQ0uMXFJQuNSTAoyAYfNuZwHwpSXSofUKHhStYUVRAYIU5L/nXa4eMNNOo7p8M1C
CbEWOdAs+4yQXIoo6q7KCmVCQbjP8PGP6mmR4nRRpQsacmP2BJz4SONhorcHYJa2t2D7BX+IQ7Sc
Nuod/8q9drOmpdRhLXjsexSLvtCx2LcfEsEQyiNPLj3X1OYUq97QO0HxVbql+QT0a52v6mT1ZW9R
AJPsX980RskhppMTnz0rp3g63nEwWV9rTQg+2jSMHWqURZMfSCZupka9Y7kmiyEs9XPVPyGwGZfl
5c88wE4WNpz0nrNU1TFTb2sL3fmeaOcr1OIYXnDXg+ONizohzVgU4aJxBggEjPRG1as0cC4DbMtx
/2R/YnhGjc3csi8BJKEmhqfs/m90KlysBGlTHnRlhFwuHGrv2sktvyqRfmrWJkPPNQx9anCHkD3x
dKrflfaA9hvT0ASTRWRK1i7fRchfho6H66oryZuwgVENja+ZXYiLFL6Q7TYrdaoLkNlJ3wapIRYo
KemmnQA40U7BBzMBRDSP/fZamYCQQC/nIdS6GhzyxHpx/vpcj1yRfpDBIIbblkSrO2CSU+Y7Tu1n
NwWg1E8yb8xaFt6jHPAbmUY/vZllhKJ6x72CF5+ek+e6dGAymJx2Q8jP35BAPHtK6XEPXUAcd439
mpWz2unTyCtfuLRXhxTUGQ4QE5EoYWv7TkaKniax6cMNG8q25fFF+LKmOWXwHzmeZ8KHh0uMFI+o
vW7aZwHNGnm3KOgVhX+Ug0Nwfgt2vgeJWPM8MbR/2mFUswl8OOoij4xHfBCA0oSeGODYOwZWr9b8
kpTsCqUEFpOR48Xlspip41ZzmOA6Tf2xcil4V07J622H+F/W/qPCt6R34xL2vAldgWCJvBiPANgJ
zQF0MOPqck9OMLasd8JOakURa5nNB2J70UyL9DcP5O/hnY+C2uSw9vNKDTVgDdofeI7bvLSrWNAO
cEyAQoqajotQhn6W5G8Zc+xnQg1/pDuwsG0Y5a/2fCs5EIgCskEOm2L7kUtzMhuNCuxk4uLnK4iX
avTbC1QlZinmYa+ULCK6LosemlFGj0lDTDlcCD8h6Lpxah0jwet6ufFPkQ6Z81PWaub1KNuYGcgH
UcZGmNwEVo4c6WnLq1XSKrxInpdXDwPi2SopvH7xr0pxnwJO7bbbGga3zRvqDtYONaP2b3paC8OI
PBj6RNkTZCCTMtscDVkF8MxeE1UQEiLqLQJCHV3Lkeb4ZK+yqbLOVcZcAzdNiltsvJxiATZaSQz2
5EzDmUsXcjxW45Kv7DIzMgFzS1f2L/RSmr4KdarWcZDNW9QBB65MGJCsfi2NDVpFlaxx+51h4uvg
qIwRxQjO0P5Sp+boyT63U3u7yY3GdldiYOUU5meknfeXLcARDudcyM4WBmT1MN5B9VZiXyMk7wUB
5Lf4iJr1NTnKekbMJkuktI0uk3lIc4GEQGKfwjBWLlvR4kojhUxbteV9zdskxbYyCEM8FHiQHdRw
bL86Ac/ksKUcUGWEOxvyWGve+YsLtIFLyNywGyHx7KP3UHj8Snq63YGWQFWBeZbaL+jnT1RK3wLP
6yA5ZqP+Ok9BZO5+EpWDeofR6JCWqIz/MiB7wsVgezKC9Vfpe4ljSCUByFjufX+B/XJE2ST2atWT
fKcw9WW3E2I33vniuIIBtYDqf5IN1EsBvr3UrtuxDgvjbMEtY0b4M0XdBl94dnq3GXEAh72sFrmw
B9lO4Wl9YhJgHfPzktuzSdmoERJES61ugf3qZ6u+UZOiVF4wBgJsrY7hAbFswWYDBPHrLUnCk1TD
CR96dn8LGBLmlGNebNkBY7aZw+uVg5hqpE7ExbicXxADFAciDE86n5Kj9maHIrINSiVHy/zBqUHY
k+UGCdRrgr7gTVjTvdc7FpiV4Pb4eFSz3P9VqW3gtw8/quXMnz307Nqzjn7rxjItu57R6FsotHTo
Ss1WQRl6nqZh/ygj0jVethRxwohKd3CXzTr9wr74zHY8XksCm3iXAJsW1dfXXxOKoiWf0IbUBxic
mYLFVOvbHr1afXQuy1EmVxI5VY+2l39YwfeY2SUTdCrJgqcOBEmTnMHD5AN2Fqa+NbkTBjxkmivE
om4l5rsCdLnVpIPmbTCWhXNwun/eZnNVvvRFnasiFJ9ekjGtMIyOAo0SnFyHTfGjmrTmsIvy/JYb
yijLdHY14eVGnM38DeQH8ibzOvSl7lp0SEQoId6VzuEen1kew9ioe0jY4ZZz8+XrOMsXPrPD4H9x
msUUBBPphVrpk4M97AvNp2lRfsAvg+7K7ZbNBJCPV5xmhFcFW/ObIyN79vYAxlTxyNT22IBdKDlU
/KOo9eOICe/u8lmv2/eRgzEh3dvoN6HK4W1GOZ2qaRhH0EsL8cYHkCS/QV1z1H393/n1+FIlpZaO
t0DhZtRdZ+AJgyMA+B2nX8B6AI2VuZIz216D8vpAW/tudwKI0Mma6E/9pwD2WwR4LK79p5lcbXcl
UAcW+i6v19IZszTkbxFKpnKPKplNnH3DyNM/Ur9zA47L22/5uy95IfU27+jx23l0uWCSmFbof81z
EuDk8mmPF3w9U33M4PvBjOLayVH1Bi2T/RQ4VJyFhwJ1nXhbxcNrFIJtU2OqQ0ddHIxYqbQtKzsD
pTuZ8//vD9ccc/gaJb74oWS+gWhU/DsrHt5pix2gK6xq9yE2JgMNF/ZHRavnQfFe6XuL+hW6vBIm
/q3/XOTwUuleLb3JrmgUBpdW0W8zA9bd4hwsZ9rXSjA/6EovibZQJFyJ5WliQmEpd7S5N/Dk5C5x
eFdq2LnlPUVzPjexNOzZzlwGqyyxPSvd0HLv33t8VoaPbU2rOwE8vyUJ1DgNl7NFgaLlNWZnGPOj
EohXmEVgIyaD4y9WdpIWPnKoTd1sNu0dgGmUlriLrlmrwzWamhQrrN2la/AOvNXLgHLzo7Li33cG
Q1xoF847pCFVIrFqsKVW8zmAgxmVfVXsv1Wmgbvkkn6vqkLhjZdc/n4yUIt1yVHi5/xqfeq+y+id
5cW16HxBBcaQ1LyXKFEL/Mlr1Z0VWUw+SwiVYGOtrw77EzdYBOZ3GDpFvfqBgoOigQtgNJ8vMbH0
uNjxoOlCr/A6QLwQ9is/yaGt0SvkQWMDJCogWvofHONTHo0DL4cfELtKzWlnEeLJYrV/XNcDigl2
eCSkKJ9ZvFJC682KgjTJOSPIr3SwdZ0lqRKd7oW1kCLvJmgr1iL0y/fhJkxFobOC1AA3HhSoYGOx
aDfYMqakuQF80dTHzBeV5oSw3+2mPpCmSRlKYcDlWqDB01y4bil7RFt+VG38/Oxf64o7GUALB/No
dIR9eG5oCuL/tZwXQHFF4hSYJ0ngW8bf/aaUZL/WjFXCiFfbWWY/eqXUImgaNKHn1AwSQSbFPnj9
bRWNL6eqax9EITE1XRRMO4MCisNDrHQM15n49cyAOraJB/q0mIfwCQlpu0SiADUiiaJmbSu2RSPM
Vz1mQCmBb5gyd5RGSxtcj/qtZYpg+6haerft9YTl0A0hhhkMi5VWQU86sWjzEbYm7gGftg0khmAa
IPaSUSjd63qamG71OMjAdIXCUX+G7zl0+oQWG0sJRnD4TjdhFE4ulzy9Wlxq8Ojo5I5k3/LfjL46
kkf79cClhIlDbkodGj8x0cXz/gdUXhZwHom6nuTazPme73xxXnMg482mbb5LgDCnaI6JDaZ8ehCe
r2JUf4Ujd9EdUfIE+EW8MxvXZC6z03lOZOuIWypbKh69NdOGiMemDfviIHJXeVbpAy8DShBnUt7t
JDXwl1CVdzgPFyXclfp/vxTLyNHLM3xHzMElukhldpovH1ffILlqjv4hyaw6xZqNs7JUh4y7PAw6
jbpqAb7G0tQCMjZfuDlo8qmPeAK8561jUKVleoc3wsYnzZGQ9pAVpmpasEuwoZVQfNXph6aMlg+G
GL7v3de/oJU/OZdpAwlkhW1Kx5vNH8Wm5gv74I3g9++pcF2cafA4KYoUCHxN3OLnpMLUdIUj0LSP
sK/PrBqj
`pragma protect end_protected

