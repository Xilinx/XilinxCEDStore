wire cpm5pldma0resetn;
wire cpm5pldma1resetn;

wire gt_refclk0_div2_ibuf;
wire gt_refclk1_div2_ibuf;

wire [11:0] cpm5rclk0;
wire [11:0] cpm5rclk1;
wire [31:0] cpm5plgpo0;
wire [31:0] cpm5plgpo1;

wire ifcpm5plaxi0wlast;
wire ifcpm5plaxi0arlock;
wire ifcpm5plaxi0awlock;
wire ifcpm5plaxi0bready;
wire ifcpm5plaxi0bvalid;
wire ifcpm5plaxi0rready;
wire ifcpm5plaxi0rvalid;
wire ifcpm5plaxi0wready;
wire ifcpm5plaxi0wvalid;
wire ifcpm5plaxi0arready;
wire ifcpm5plaxi0arvalid;
wire ifcpm5plaxi0awready;
wire ifcpm5plaxi0awvalid;
wire [15:0] ifcpm5plaxi0bid;
wire [15:0] ifcpm5plaxi0rid;
wire [15:0] ifcpm5plaxi0wid;
wire [15:0] ifcpm5plaxi0arid;
wire [15:0] ifcpm5plaxi0awid;
wire [0:0]  ifcpm5plaxi0buser;
wire [0:0]  ifcpm5plaxi0rlast;
wire [1:0]  ifcpm5plaxi0bresp;
wire [1:0]  ifcpm5plaxi0rresp;
wire [3:0]  ifcpm5plaxi0arqos;
wire [3:0]  ifcpm5plaxi0awqos;
wire [63:0] ifcpm5plaxi0wstrb;
wire [7:0]  ifcpm5plaxi0arlen;
wire [7:0]  ifcpm5plaxi0awlen;
wire[127:0] ifcpm5plaxi0ruser;
wire[127:0] ifcpm5plaxi0wuser;
wire[511:0] ifcpm5plaxi0rdata;
wire[511:0] ifcpm5plaxi0wdata;
wire [2:0]  ifcpm5plaxi0arprot;
wire [2:0]  ifcpm5plaxi0arsize;
wire [2:0]  ifcpm5plaxi0awprot;
wire [2:0]  ifcpm5plaxi0awsize;
wire [31:0] ifcpm5plaxi0aruser;
wire [31:0] ifcpm5plaxi0awuser;
wire [63:0] ifcpm5plaxi0araddr;
wire [63:0] ifcpm5plaxi0awaddr;
wire [1:0]  ifcpm5plaxi0arburst;
wire [1:0]  ifcpm5plaxi0awburst;
wire [3:0]  ifcpm5plaxi0arcache;
wire [3:0]  ifcpm5plaxi0awcache;
wire [3:0]  ifcpm5plaxi0arregion;
wire [3:0]  ifcpm5plaxi0awregion;

wire ifcpm5plaxi1buser;
wire ifcpm5plaxi1rlast;
wire ifcpm5plaxi1bready;
wire ifcpm5plaxi1bvalid;
wire ifcpm5plaxi1rready;
wire ifcpm5plaxi1rvalid;
wire ifcpm5plaxi1wready;
wire ifcpm5plaxi1wvalid;
wire ifcpm5plaxi1arready;
wire ifcpm5plaxi1arvalid;
wire ifcpm5plaxi1awready;
wire ifcpm5plaxi1awvalid;
wire [15:0] ifcpm5plaxi1bid;
wire [15:0] ifcpm5plaxi1rid;
wire [15:0] ifcpm5plaxi1wid;
wire [15:0] ifcpm5plaxi1arid;
wire [15:0] ifcpm5plaxi1awid;
wire [0:0]  ifcpm5plaxi1wlast;
wire [1:0]  ifcpm5plaxi1bresp;
wire [1:0]  ifcpm5plaxi1rresp;
wire [3:0]  ifcpm5plaxi1arqos;
wire [3:0]  ifcpm5plaxi1awqos;
wire [63:0] ifcpm5plaxi1wstrb;
wire [7:0]  ifcpm5plaxi1arlen;
wire [7:0]  ifcpm5plaxi1awlen;
wire[127:0] ifcpm5plaxi1ruser;
wire[127:0] ifcpm5plaxi1wuser;
wire[511:0] ifcpm5plaxi1rdata;
wire[511:0] ifcpm5plaxi1wdata;
wire [0:0]  ifcpm5plaxi1arlock;
wire [0:0]  ifcpm5plaxi1awlock;
wire [2:0]  ifcpm5plaxi1arprot;
wire [2:0]  ifcpm5plaxi1arsize;
wire [2:0]  ifcpm5plaxi1awprot;
wire [2:0]  ifcpm5plaxi1awsize;
wire [31:0] ifcpm5plaxi1aruser;
wire [31:0] ifcpm5plaxi1awuser;
wire [63:0] ifcpm5plaxi1araddr;
wire [63:0] ifcpm5plaxi1awaddr;
wire [1:0]  ifcpm5plaxi1arburst;
wire [1:0]  ifcpm5plaxi1awburst;
wire [3:0]  ifcpm5plaxi1arcache;
wire [3:0]  ifcpm5plaxi1awcache;
wire [3:0]  ifcpm5plaxi1arregion;
wire [3:0]  ifcpm5plaxi1awregion;

wire ifcpm5plisrcorrevent;
wire ifcpm5plisrmiscevent;
wire ifcpm5plisruncorrevent;

wire ifcpm5plmpio0cfgfcvcsel;
wire ifcpm5plmpio0cfgflrdone;
wire ifcpm5plmpio0axiscctlast;
wire ifcpm5plmpio0axiscqtlast;
wire ifcpm5plmpio0axisrctlast;
wire ifcpm5plmpio0axisrqtlast;
wire ifcpm5plmpio0cfgerrcorin;
wire ifcpm5plmpio0cfgmgmtread;
wire ifcpm5plmpio0cfgreqrxack;
wire ifcpm5plmpio0axiscctvalid;
wire ifcpm5plmpio0axisrqtvalid;
wire ifcpm5plmpio0cfgedrenable;
wire ifcpm5plmpio0cfgerrcorout;
wire ifcpm5plmpio0cfgmgmt2read;
wire ifcpm5plmpio0cfgmgmtwrite;
wire ifcpm5plmpio0cfgrcbstatus;
wire ifcpm5plmpio0cfgvc1enable;
wire ifcpm5plmpio0cfgerruncorin;
wire ifcpm5plmpio0cfghotresetin;
wire ifcpm5plmpio0cfgmgmt2write;
wire ifcpm5plmpio0cfgperfuncreq;
wire ifcpm5plmpio0cfgperfuncvld;
wire ifcpm5plmpio0pcieaxiscqrts;
wire ifcpm5plmpio0pcieaxiscqvld;
wire ifcpm5plmpio0pcieaxisrcrts;
wire ifcpm5plmpio0pcieaxisrcvld;
wire ifcpm5plmpio0cfgerrfatalout;
wire ifcpm5plmpio0cfghotresetout;
wire ifcpm5plmpio0cfgmsgreceived;
wire ifcpm5plmpio0cfgmsgtransmit;
wire ifcpm5plmpio0cfgpasidenable;
wire ifcpm5plmpio0cfgphylinkdown;
wire ifcpm5plmpio0cfgreqrxtready;
wire ifcpm5plmpio0cfgreqrxtvalid;
wire ifcpm5plmpio0cfgreqtxtready;
wire ifcpm5plmpio0cfgreqtxtvalid;
wire ifcpm5plmpio0cfgwrreqbmevld;
wire ifcpm5plmpio0cfgwrreqflrvld;
wire ifcpm5plmpio0cfgwrreqmsivld;
wire ifcpm5plmpio0cfgwrreqvfevld;
wire ifcpm5plmpio0cfgexttagenable;
wire ifcpm5plmpio0cfgwrreqmsixvld;
wire ifcpm5plmpio0cfgerrmsgtypevld;
wire ifcpm5plmpio0cfginterruptsent;
wire ifcpm5plmpio0cfgerrnonfatalout;
wire ifcpm5plmpio0cfgplstatuschange;
wire ifcpm5plmpio0cfgextreadreceived;
wire ifcpm5plmpio0cfglocalerrorvalid;
wire ifcpm5plmpio0cfgmgmtdebugaccess;
wire ifcpm5plmpio0cfgmsgtransmitdone;
wire ifcpm5plmpio0cfgextreaddatavalid;
wire ifcpm5plmpio0cfgextwritereceived;
wire ifcpm5plmpio0cfginterruptmsifail;
wire ifcpm5plmpio0cfginterruptmsisent;
wire ifcpm5plmpio0cfginterruptmsixint;
wire ifcpm5plmpio0cfgmgmt2debugaccess;
wire ifcpm5plmpio0cfginterruptmsixmask;
wire ifcpm5plmpio0cfgmgmtreadwritedone;
wire ifcpm5plmpio0cfginterruptmsienable;
wire ifcpm5plmpio0cfgmgmt2readwritedone;
wire ifcpm5plmpio0cfginterruptmsixenable;
wire ifcpm5plmpio0cfgpowerstatechangeack;
wire ifcpm5plmpio0cfg10btagrequesterenable;
wire ifcpm5plmpio0cfgatomicrequesterenable;
wire ifcpm5plmpio0cfgpasidprivilmodeenable;
wire ifcpm5plmpio0cfgvc1negotiationpending;
wire ifcpm5plmpio0cfginterruptmsimaskupdate;
wire ifcpm5plmpio0cfginterruptmsitphpresent;
wire ifcpm5plmpio0cfgccixedrdataratechangeack;
wire ifcpm5plmpio0cfgccixedrdataratechangereq;
wire ifcpm5plmpio0cfgpasidexecpermissionenable;
wire ifcpm5plmpio0cfgpowerstatechangeinterrupt;
wire ifcpm5plmpio0cfginterruptmsixvecpendingstatus;
wire ifcpm5plmpio0cfginterruptmsipendingstatusdataenable;

wire [11:0]  ifcpm5plmpio0cfgfcpd;
wire [7:0]   ifcpm5plmpio0cfgfcph;
wire [11:0]  ifcpm5plmpio0cfgfcnpd;
wire [2:0]   ifcpm5plmpio0cfgfcsel;
wire [7:0]   ifcpm5plmpio0cfgfcnph;
wire [11:0]  ifcpm5plmpio0cfgfccpld;
wire [39:0]  ifcpm5plmpio0pcierqtag;
wire [7:0]   ifcpm5plmpio0cfgfccplh;
wire [164:0] ifcpm5plmpio0axiscctuser;
wire [2:0]   ifcpm5plmpio0pciecqnpreq;
wire [3:0]   ifcpm5plmpio0pcierqtagav;
wire [31:0]  ifcpm5plmpio0axiscctkeep;
wire [31:0]  ifcpm5plmpio0axiscqtkeep;
wire [31:0]  ifcpm5plmpio0axisrqtkeep;
wire [372:0] ifcpm5plmpio0axisrqtuser;
wire [9:0]   ifcpm5plmpio0cfgmgmtaddr;
wire[1023:0] ifcpm5plmpio0axiscctdata;
wire[1023:0] ifcpm5plmpio0axiscqtdata;
wire[1023:0] ifcpm5plmpio0axisrqtdata;
wire[464:0]  ifcpm5plmpio0axiscqtuser;
wire [1:0]   ifcpm5plmpio0cfgfcpdscale;
wire [1:0]   ifcpm5plmpio0cfgfcphscale;
wire [1:0]   ifcpm5plmpio0cfgrxpmstate;
wire [1:0]   ifcpm5plmpio0cfgtxpmstate;
wire [3:0]   ifcpm5plmpio0pcierqtagvld;
wire [3:0]   ifcpm5plmpio0pcietfcnpdav;
wire [3:0]   ifcpm5plmpio0pcietfcnphav;
wire [7:0]   ifcpm5plmpio0axiscctready;
wire [7:0]   ifcpm5plmpio0axisrqtready;
wire [7:0]   ifcpm5plmpio0cfgbusnumber;
wire [9:0]   ifcpm5plmpio0cfgmgmt2addr;
wire [1:0]   ifcpm5plmpio0cfgfcnpdscale;
wire [1:0]   ifcpm5plmpio0cfgfcnphscale;
wire [1:0]   ifcpm5plmpio0cfgmaxpayload;
wire [127:0] ifcpm5plmpio0cfgreqrxtdata;
wire [127:0] ifcpm5plmpio0cfgreqtxtdata;
wire [16:0]  ifcpm5plmpio0cfgreqrxtuser;
wire [16:0]  ifcpm5plmpio0cfgreqtxtuser;
wire [2:0]   ifcpm5plmpio0cfgmaxreadreq;
wire [23:0]  ifcpm5plmpio0cfgperfuncout;
wire [5:0]   ifcpm5plmpio0cfgerrmsgtype;
wire [5:0]   ifcpm5plmpio0cfgltssmstate;
wire [5:0]   ifcpm5plmpio0pcierqseqnum0;
wire [5:0]   ifcpm5plmpio0pcierqseqnum1;
wire [5:0]   ifcpm5plmpio0pcierqseqnum2;
wire [5:0]   ifcpm5plmpio0pcierqseqnum3;
wire [1:0]   ifcpm5plmpio0cfgfccpldscale;
wire [1:0]   ifcpm5plmpio0cfgfccplhscale;
wire [31:0]  ifcpm5plmpio0cfgextreaddata;
wire [15:0]  ifcpm5plmpio0cfgwrreqfuncnum;
wire [2:0]   ifcpm5plmpio0cfgcurrentspeed;
wire [3:0]   ifcpm5plmpio0cfginterruptint;
wire [3:0]   ifcpm5plmpio0pcierqseqnumvld;
wire [31:0]  ifcpm5plmpio0cfgextwritedata;
wire [31:0]  ifcpm5plmpio0cfgmgmtreaddata;
wire [59:0]  ifcpm5plmpio0pcieaxiscqready;
wire [59:0]  ifcpm5plmpio0pcieaxisrcready;
wire [1:0]   ifcpm5plmpio0cfgphylinkstatus;
wire [3:0]   ifcpm5plmpio0cfgwrreqoutvalue;
wire [31:0]  ifcpm5plmpio0cfgmgmt2readdata;
wire [31:0]  ifcpm5plmpio0cfgmgmtwritedata;
wire [4:0]   ifcpm5plmpio0cfglocalerrorout;
wire [5:0]   ifcpm5plmpio0pciecqnpreqcount;
wire [1:0]   ifcpm5plmpio0cfglinkpowerstate;
wire [15:0]  ifcpm5plmpio0cfgflrdonefuncnum;
wire [15:0]  ifcpm5plmpio0cfgperfuncfuncnum;
wire [3:0]   ifcpm5plmpio0cfgfunctionstatus;
wire [3:0]   ifcpm5plmpio0cfgmgmtbyteenable;
wire [31:0]  ifcpm5plmpio0cfgmgmt2writedata;
wire [2:0]   ifcpm5plmpio0cfgmsgtransmittype;
wire [2:0]   ifcpm5plmpio0cfgnegotiatedwidth;
wire [3:0]   ifcpm5plmpio0cfgmgmt2byteenable;
wire [31:0]  ifcpm5plmpio0cfginterruptmsiint;
wire [31:0]  ifcpm5plmpio0cfgmsgtransmitdata;
wire [4:0]   ifcpm5plmpio0cfgmsgreceivedtype;
wire [7:0]   ifcpm5plmpio0cfgmsgreceiveddata;
wire [15:0]  ifcpm5plmpio0cfginterruptpending;
wire [2:0]   ifcpm5plmpio0cfginterruptmsiattr;
wire [31:0]  ifcpm5plmpio0cfginterruptmsidata;
wire [15:0]  ifcpm5plmpio0cfgextfunctionnumber;
wire [31:0]  ifcpm5plmpio0cfginterruptmsixdata;
wire [9:0]   ifcpm5plmpio0cfgextregisternumber;
wire [15:0]  ifcpm5plmpio0cfgmgmtfunctionnumber;
wire [2:0]   ifcpm5plmpio0cfgfunctionpowerstate;
wire [3:0]   ifcpm5plmpio0cfgextwritebyteenable;
wire [3:0]   ifcpm5plmpio0cfginterruptmsiselect;
wire [1:0]   ifcpm5plmpio0cfginterruptmsitphtype;
wire [15:0]  ifcpm5plmpio0cfgmgmt2functionnumber;
wire [2:0]   ifcpm5plmpio0cfginterruptmsimmenable;
wire [63:0]  ifcpm5plmpio0cfginterruptmsixaddress;
wire [7:0]   ifcpm5plmpio0cfginterruptmsitphsttag;
wire [9:0]   ifcpm5plmpio0cfgerrmsgfunctionnumber;
wire [1:0]   ifcpm5plmpio0cfginterruptmsixvecpending;
wire [31:0]  ifcpm5plmpio0cfginterruptmsipendingstatus;
wire [15:0]  ifcpm5plmpio0cfginterruptmsifunctionnumber;
wire [3:0]   ifcpm5plmpio0cfginterruptmsipendingstatusfunctionnum;

wire ifcpm5plmpio1cfgfcvcsel;
wire ifcpm5plmpio1cfgflrdone;
wire ifcpm5plmpio1axiscctlast;
wire ifcpm5plmpio1axiscqtlast;
wire ifcpm5plmpio1axisrctlast;
wire ifcpm5plmpio1axisrqtlast;
wire ifcpm5plmpio1cfgerrcorin;
wire ifcpm5plmpio1cfgmgmtread;
wire ifcpm5plmpio1cfgreqrxack;
wire ifcpm5plmpio1axiscctvalid;
wire ifcpm5plmpio1axisrqtvalid;
wire ifcpm5plmpio1cfgedrenable;
wire ifcpm5plmpio1cfgerrcorout;
wire ifcpm5plmpio1cfgmgmt2read;
wire ifcpm5plmpio1cfgmgmtwrite;
wire ifcpm5plmpio1cfgrcbstatus;
wire ifcpm5plmpio1cfgvc1enable;
wire ifcpm5plmpio1cfgerruncorin;
wire ifcpm5plmpio1cfghotresetin;
wire ifcpm5plmpio1cfgmgmt2write;
wire ifcpm5plmpio1cfgperfuncreq;
wire ifcpm5plmpio1cfgperfuncvld;
wire ifcpm5plmpio1pcieaxiscqrts;
wire ifcpm5plmpio1pcieaxiscqvld;
wire ifcpm5plmpio1pcieaxisrcrts;
wire ifcpm5plmpio1pcieaxisrcvld;
wire ifcpm5plmpio1cfgerrfatalout;
wire ifcpm5plmpio1cfghotresetout;
wire ifcpm5plmpio1cfgmsgreceived;
wire ifcpm5plmpio1cfgmsgtransmit;
wire ifcpm5plmpio1cfgpasidenable;
wire ifcpm5plmpio1cfgphylinkdown;
wire ifcpm5plmpio1cfgreqrxtready;
wire ifcpm5plmpio1cfgreqrxtvalid;
wire ifcpm5plmpio1cfgreqtxtready;
wire ifcpm5plmpio1cfgreqtxtvalid;
wire ifcpm5plmpio1cfgwrreqbmevld;
wire ifcpm5plmpio1cfgwrreqflrvld;
wire ifcpm5plmpio1cfgwrreqmsivld;
wire ifcpm5plmpio1cfgwrreqvfevld;
wire ifcpm5plmpio1cfgexttagenable;
wire ifcpm5plmpio1cfgwrreqmsixvld;
wire ifcpm5plmpio1cfgerrmsgtypevld;
wire ifcpm5plmpio1cfginterruptsent;
wire ifcpm5plmpio1cfgerrnonfatalout;
wire ifcpm5plmpio1cfgplstatuschange;
wire ifcpm5plmpio1cfgextreadreceived;
wire ifcpm5plmpio1cfglocalerrorvalid;
wire ifcpm5plmpio1cfgmgmtdebugaccess;
wire ifcpm5plmpio1cfgmsgtransmitdone;
wire ifcpm5plmpio1cfgextreaddatavalid;
wire ifcpm5plmpio1cfgextwritereceived;
wire ifcpm5plmpio1cfginterruptmsifail;
wire ifcpm5plmpio1cfginterruptmsisent;
wire ifcpm5plmpio1cfginterruptmsixint;
wire ifcpm5plmpio1cfgmgmt2debugaccess;
wire ifcpm5plmpio1cfginterruptmsixmask;
wire ifcpm5plmpio1cfgmgmtreadwritedone;
wire ifcpm5plmpio1cfginterruptmsienable;
wire ifcpm5plmpio1cfgmgmt2readwritedone;
wire ifcpm5plmpio1cfginterruptmsixenable;
wire ifcpm5plmpio1cfgpowerstatechangeack;
wire ifcpm5plmpio1cfg10btagrequesterenable;
wire ifcpm5plmpio1cfgatomicrequesterenable;
wire ifcpm5plmpio1cfgpasidprivilmodeenable;
wire ifcpm5plmpio1cfgvc1negotiationpending;
wire ifcpm5plmpio1cfginterruptmsimaskupdate;
wire ifcpm5plmpio1cfginterruptmsitphpresent;
wire ifcpm5plmpio1cfgccixedrdataratechangeack;
wire ifcpm5plmpio1cfgccixedrdataratechangereq;
wire ifcpm5plmpio1cfgpasidexecpermissionenable;
wire ifcpm5plmpio1cfgpowerstatechangeinterrupt;
wire ifcpm5plmpio1cfginterruptmsixvecpendingstatus;
wire ifcpm5plmpio1cfginterruptmsipendingstatusdataenable;

wire [11:0]  ifcpm5plmpio1cfgfcpd;
wire [7:0]   ifcpm5plmpio1cfgfcph;
wire [11:0]  ifcpm5plmpio1cfgfcnpd;
wire [2:0]   ifcpm5plmpio1cfgfcsel;
wire [7:0]   ifcpm5plmpio1cfgfcnph;
wire [11:0]  ifcpm5plmpio1cfgfccpld;
wire [39:0]  ifcpm5plmpio1pcierqtag;
wire [7:0]   ifcpm5plmpio1cfgfccplh;
wire [164:0] ifcpm5plmpio1axiscctuser;
wire [2:0]   ifcpm5plmpio1pciecqnpreq;
wire [3:0]   ifcpm5plmpio1pcierqtagav;
wire [31:0]  ifcpm5plmpio1axiscctkeep;
wire [31:0]  ifcpm5plmpio1axiscqtkeep;
wire [31:0]  ifcpm5plmpio1axisrqtkeep;
wire [372:0] ifcpm5plmpio1axisrqtuser;
wire [9:0]   ifcpm5plmpio1cfgmgmtaddr;
wire[1023:0] ifcpm5plmpio1axiscctdata;
wire[1023:0] ifcpm5plmpio1axiscqtdata;
wire[1023:0] ifcpm5plmpio1axisrqtdata;
wire[464:0]  ifcpm5plmpio1axiscqtuser;
wire [1:0]   ifcpm5plmpio1cfgfcpdscale;
wire [1:0]   ifcpm5plmpio1cfgfcphscale;
wire [1:0]   ifcpm5plmpio1cfgrxpmstate;
wire [1:0]   ifcpm5plmpio1cfgtxpmstate;
wire [3:0]   ifcpm5plmpio1pcierqtagvld;
wire [3:0]   ifcpm5plmpio1pcietfcnpdav;
wire [3:0]   ifcpm5plmpio1pcietfcnphav;
wire [7:0]   ifcpm5plmpio1axiscctready;
wire [7:0]   ifcpm5plmpio1axisrqtready;
wire [7:0]   ifcpm5plmpio1cfgbusnumber;
wire [9:0]   ifcpm5plmpio1cfgmgmt2addr;
wire [1:0]   ifcpm5plmpio1cfgfcnpdscale;
wire [1:0]   ifcpm5plmpio1cfgfcnphscale;
wire [1:0]   ifcpm5plmpio1cfgmaxpayload;
wire [127:0] ifcpm5plmpio1cfgreqtxtdata;
wire [16:0]  ifcpm5plmpio1cfgreqrxtuser;
wire [16:0]  ifcpm5plmpio1cfgreqtxtuser;
wire [2:0]   ifcpm5plmpio1cfgmaxreadreq;
wire [23:0]  ifcpm5plmpio1cfgperfuncout;
wire [5:0]   ifcpm5plmpio1cfgerrmsgtype;
wire [5:0]   ifcpm5plmpio1cfgltssmstate;
wire [5:0]   ifcpm5plmpio1pcierqseqnum0;
wire [5:0]   ifcpm5plmpio1pcierqseqnum1;
wire [5:0]   ifcpm5plmpio1pcierqseqnum2;
wire [5:0]   ifcpm5plmpio1pcierqseqnum3;
wire [127:0] ifcpm5plmpio1cfgreqrxtdata;
wire [1:0]   ifcpm5plmpio1cfgfccpldscale;
wire [1:0]   ifcpm5plmpio1cfgfccplhscale;
wire [31:0]  ifcpm5plmpio1cfgextreaddata;
wire [15:0]  ifcpm5plmpio1cfgwrreqfuncnum;
wire [2:0]   ifcpm5plmpio1cfgcurrentspeed;
wire [3:0]   ifcpm5plmpio1cfginterruptint;
wire [3:0]   ifcpm5plmpio1pcierqseqnumvld;
wire [31:0]  ifcpm5plmpio1cfgextwritedata;
wire [31:0]  ifcpm5plmpio1cfgmgmtreaddata;
wire [59:0]  ifcpm5plmpio1pcieaxiscqready;
wire [59:0]  ifcpm5plmpio1pcieaxisrcready;
wire [1:0]   ifcpm5plmpio1cfgphylinkstatus;
wire [3:0]   ifcpm5plmpio1cfgwrreqoutvalue;
wire [31:0]  ifcpm5plmpio1cfgmgmt2readdata;
wire [31:0]  ifcpm5plmpio1cfgmgmtwritedata;
wire [4:0]   ifcpm5plmpio1cfglocalerrorout;
wire [5:0]   ifcpm5plmpio1pciecqnpreqcount;
wire [1:0]   ifcpm5plmpio1cfglinkpowerstate;
wire [15:0]  ifcpm5plmpio1cfgflrdonefuncnum;
wire [15:0]  ifcpm5plmpio1cfgperfuncfuncnum;
wire [3:0]   ifcpm5plmpio1cfgfunctionstatus;
wire [3:0]   ifcpm5plmpio1cfgmgmtbyteenable;
wire [31:0]  ifcpm5plmpio1cfgmgmt2writedata;
wire [2:0]   ifcpm5plmpio1cfgmsgtransmittype;
wire [2:0]   ifcpm5plmpio1cfgnegotiatedwidth;
wire [3:0]   ifcpm5plmpio1cfgmgmt2byteenable;
wire [31:0]  ifcpm5plmpio1cfginterruptmsiint;
wire [31:0]  ifcpm5plmpio1cfgmsgtransmitdata;
wire [4:0]   ifcpm5plmpio1cfgmsgreceivedtype;
wire [7:0]   ifcpm5plmpio1cfgmsgreceiveddata;
wire [15:0]  ifcpm5plmpio1cfginterruptpending;
wire [2:0]   ifcpm5plmpio1cfginterruptmsiattr;
wire [31:0]  ifcpm5plmpio1cfginterruptmsidata;
wire [15:0]  ifcpm5plmpio1cfgextfunctionnumber;
wire [31:0]  ifcpm5plmpio1cfginterruptmsixdata;
wire [9:0]   ifcpm5plmpio1cfgextregisternumber;
wire [15:0]  ifcpm5plmpio1cfgmgmtfunctionnumber;
wire [2:0]   ifcpm5plmpio1cfgfunctionpowerstate;
wire [3:0]   ifcpm5plmpio1cfgextwritebyteenable;
wire [3:0]   ifcpm5plmpio1cfginterruptmsiselect;
wire [1:0]   ifcpm5plmpio1cfginterruptmsitphtype;
wire [15:0]  ifcpm5plmpio1cfgmgmt2functionnumber;
wire [2:0]   ifcpm5plmpio1cfginterruptmsimmenable;
wire [63:0]  ifcpm5plmpio1cfginterruptmsixaddress;
wire [7:0]   ifcpm5plmpio1cfginterruptmsitphsttag;
wire [9:0]   ifcpm5plmpio1cfgerrmsgfunctionnumber;
wire [1:0]   ifcpm5plmpio1cfginterruptmsixvecpending;
wire [31:0]  ifcpm5plmpio1cfginterruptmsipendingstatus;
wire [15:0]  ifcpm5plmpio1cfginterruptmsifunctionnumber;
wire [3:0]   ifcpm5plmpio1cfginterruptmsipendingstatusfunctionnum;

wire ifcpmpsaxi0buser;
wire ifcpmpsaxi0rlast;
wire ifcpmpsaxi0bready;
wire ifcpmpsaxi0bvalid;
wire ifcpmpsaxi0rready;
wire ifcpmpsaxi0rvalid;
wire ifcpmpsaxi0wready;
wire ifcpmpsaxi0wvalid;
wire ifcpmpsaxi0arready;
wire ifcpmpsaxi0arvalid;
wire ifcpmpsaxi0awready;
wire ifcpmpsaxi0awvalid;
wire [15:0] ifcpmpsaxi0bid;
wire [15:0] ifcpmpsaxi0rid;
wire [15:0] ifcpmpsaxi0wid;
wire [15:0] ifcpmpsaxi0arid;
wire [15:0] ifcpmpsaxi0awid;
wire [0:0]  ifcpmpsaxi0wlast;
wire [1:0]  ifcpmpsaxi0bresp;
wire [1:0]  ifcpmpsaxi0rresp;
wire [15:0] ifcpmpsaxi0wstrb;
wire [17:0] ifcpmpsaxi0ruser;
wire [17:0] ifcpmpsaxi0wuser;
wire [3:0]  ifcpmpsaxi0arqos;
wire [3:0]  ifcpmpsaxi0awqos;
wire [7:0]  ifcpmpsaxi0arlen;
wire [7:0]  ifcpmpsaxi0awlen;
wire[127:0] ifcpmpsaxi0rdata;
wire[127:0] ifcpmpsaxi0wdata;
wire [0:0]  ifcpmpsaxi0arlock;
wire [0:0]  ifcpmpsaxi0awlock;
wire [2:0]  ifcpmpsaxi0arprot;
wire [2:0]  ifcpmpsaxi0arsize;
wire [2:0]  ifcpmpsaxi0awprot;
wire [2:0]  ifcpmpsaxi0awsize;
wire [31:0] ifcpmpsaxi0aruser;
wire [31:0] ifcpmpsaxi0awuser;
wire [63:0] ifcpmpsaxi0araddr;
wire [63:0] ifcpmpsaxi0awaddr;
wire [1:0]  ifcpmpsaxi0arburst;
wire [1:0]  ifcpmpsaxi0awburst;
wire [3:0]  ifcpmpsaxi0arcache;
wire [3:0]  ifcpmpsaxi0awcache;
wire [3:0]  ifcpmpsaxi0arregion;
wire [3:0]  ifcpmpsaxi0awregion;

wire ifcpmpsaxi1rlast;
wire ifcpmpsaxi1bready;
wire ifcpmpsaxi1bvalid;
wire ifcpmpsaxi1rready;
wire ifcpmpsaxi1rvalid;
wire ifcpmpsaxi1wready;
wire ifcpmpsaxi1wvalid;
wire ifcpmpsaxi1arready;
wire ifcpmpsaxi1arvalid;
wire ifcpmpsaxi1awready;
wire ifcpmpsaxi1awvalid;
wire [15:0] ifcpmpsaxi1bid;
wire [15:0] ifcpmpsaxi1rid;
wire [15:0] ifcpmpsaxi1wid;
wire [15:0] ifcpmpsaxi1arid;
wire [15:0] ifcpmpsaxi1awid;
wire [0:0]  ifcpmpsaxi1wlast;
wire [1:0]  ifcpmpsaxi1bresp;
wire [1:0]  ifcpmpsaxi1rresp;
wire [15:0] ifcpmpsaxi1buser;
wire [15:0] ifcpmpsaxi1wstrb;
wire [16:0] ifcpmpsaxi1ruser;
wire [16:0] ifcpmpsaxi1wuser;
wire [3:0]  ifcpmpsaxi1arqos;
wire [3:0]  ifcpmpsaxi1awqos;
wire [7:0]  ifcpmpsaxi1arlen;
wire [7:0]  ifcpmpsaxi1awlen;
wire[127:0] ifcpmpsaxi1rdata;
wire[127:0] ifcpmpsaxi1wdata;
wire [0:0]  ifcpmpsaxi1arlock;
wire [0:0]  ifcpmpsaxi1awlock;
wire [17:0] ifcpmpsaxi1aruser;
wire [17:0] ifcpmpsaxi1awuser;
wire [2:0]  ifcpmpsaxi1arprot;
wire [2:0]  ifcpmpsaxi1arsize;
wire [2:0]  ifcpmpsaxi1awprot;
wire [2:0]  ifcpmpsaxi1awsize;
wire [63:0] ifcpmpsaxi1araddr;
wire [63:0] ifcpmpsaxi1awaddr;
wire [1:0]  ifcpmpsaxi1arburst;
wire [1:0]  ifcpmpsaxi1awburst;
wire [3:0]  ifcpmpsaxi1arcache;
wire [3:0]  ifcpmpsaxi1awcache;
wire [3:0]  ifcpmpsaxi1arregion;
wire [3:0]  ifcpmpsaxi1awregion;

wire ifcpmpsisrcorrevent;
wire ifcpmpsisrmiscevent;
wire ifcpmpsisruncorrevent;

wire iffcq00enppm;
wire iffcq00perstb;
wire iffcq00bufgtce;
wire iffcq00cdrhold;
wire iffcq00cdrlock;
wire iffcq00dmonclk;
wire iffcq00rxlpmen;
wire iffcq00rxpkdet;
wire iffcq00rxqpien;
wire iffcq00rxslide;
wire iffcq00rxvalid;
wire iffcq00tstclk0;
wire iffcq00tstclk1;
wire iffcq00txswing;
wire iffcq00bufgtrst;
wire iffcq00cdrovren;
wire iffcq00cfokdone;
wire iffcq00iloreset;
wire iffcq00phyready;
wire iffcq00rxlatclk;
wire iffcq00rxusrclk;
wire iffcq00rxusrrdy;
wire iffcq00txcomsas;
wire iffcq00txlatclk;
wire iffcq00txusrclk;
wire iffcq00txusrrdy;
wire iffcq00bsrserial;
wire iffcq00cdrfreqos;
wire iffcq00cdrstepsq;
wire iffcq00cdrstepsx;
wire iffcq00comsasdet;
wire iffcq00gtrxreset;
wire iffcq00gttxreset;
wire iffcq00phystatus;
wire iffcq00rxprbserr;
wire iffcq00rxqpisenn;
wire iffcq00rxqpisenp;
wire iffcq00txcominit;
wire iffcq00txcomwake;
wire iffcq00txdccdone;
wire iffcq00txinhibit;
wire iffcq00txqpisenn;
wire iffcq00txqpisenp;
wire iffcq00aptexthold;
wire iffcq00cdrbmcdreq;
wire iffcq00cdrphreset;
wire iffcq00cdrstepdir;
wire iffcq00cominitdet;
wire iffcq00comwakedet;
wire iffcq00rxcommadet;
wire iffcq00rxelecidle;
wire iffcq00rxoobreset;
wire iffcq00rxpolarity;
wire iffcq00rxsliderdy;
wire iffcq00rxslipdone;
wire iffcq00rxsyncdone;
wire iffcq00txelecidle;
wire iffcq00txpolarity;
wire iffcq00txserpwrdn;
wire iffcq00txsyncdone;
wire iffcq00aptoverwren;
wire iffcq00cdrincpctrl;
wire iffcq00ckpinrsrvd0;
wire iffcq00ckpinrsrvd1;
wire iffcq00cssdstopclk;
wire iffcq00rxcdrphdone;
wire iffcq00rxdapireset;
wire iffcq00rxoutpcsclk;
wire iffcq00rxresetdone;
wire iffcq00rxsyncallin;
wire iffcq00txcomfinish;
wire iffcq00txdapireset;
wire iffcq00txoneszeros;
wire iffcq00txoutpcsclk;
wire iffcq00txqpibiasen;
wire iffcq00txqpiweakpu;
wire iffcq00txresetdone;
wire iffcq00txsyncallin;
wire iffcq00eyescanreset;
wire iffcq00hsdppcsreset;
wire iffcq00iloresetdone;
wire iffcq00iloresetmask;
wire iffcq00rxeqtraining;
wire iffcq00rxphdlyreset;
wire iffcq00rxprbslocked;
wire iffcq00txphdlyreset;
wire iffcq00dmonfiforeset;
wire iffcq00rxbyterealign;
wire iffcq00rxchanbondseq;
wire iffcq00rxchanrealign;
wire iffcq00rxchisaligned;
wire iffcq00rxgearboxslip;
wire iffcq00rxmldchainreq;
wire iffcq00rxtermination;
wire iffcq00txmldchainreq;
wire iffcq00txswingoutlow;
wire iffcq00eyescantrigger;
wire iffcq00resetexception;
wire iffcq00rxmldchaindone;
wire iffcq00rxphasealignpd;
wire iffcq00rxpmaresetdone;
wire iffcq00rxprbscntreset;
wire iffcq00rxprogdivreset;
wire iffcq00tcoclkfsmfrout;
wire iffcq00txchicooutrsvd;
wire iffcq00txmldchaindone;
wire iffcq00txpcsresetmask;
wire iffcq00txphasealignpd;
wire iffcq00txpmaresetdone;
wire iffcq00txprbsforceerr;
wire iffcq00txprogdivreset;
wire iffcq00txswingouthigh;
wire iffcq00rxbyteisaligned;
wire iffcq00rxdapicodereset;
wire iffcq00rxdapiresetdone;
wire iffcq00rxdelayalignerr;
wire iffcq00rxdelayalignreq;
wire iffcq00rxfinealigndone;
wire iffcq00rxphasealignerr;
wire iffcq00rxphasealignreq;
wire iffcq00txdapicodereset;
wire iffcq00txdapiresetdone;
wire iffcq00txdelayalignerr;
wire iffcq00txdelayalignreq;
wire iffcq00txphasealignerr;
wire iffcq00txphasealignreq;
wire iffcq00txtxpicodereset;
wire iffcq00eyescandataerror;
wire iffcq00rxdapicodeovrden;
wire iffcq00rxmlfinealignreq;
wire iffcq00rxphasealigndone;
wire iffcq00txdapicodeovrden;
wire iffcq00txphasealigndone;
wire iffcq00txtxpicodeovrden;
wire iffcq00xpipe5pipelineen;
wire iffcq00rxphasesetinitreq;
wire iffcq00txpausedelayalign;
wire iffcq00txphasesetinitreq;
wire iffcq00rxphasesetinitdone;
wire iffcq00rxphaseshift180req;
wire iffcq00rxprogdivresetdone;
wire iffcq00rxsimplexphystatus;
wire iffcq00txdetectrxloopback;
wire iffcq00txphasesetinitdone;
wire iffcq00txphaseshift180req;
wire iffcq00txprogdivresetdone;
wire iffcq00txsimplexphystatus;
wire iffcq00rxphaseshift180done;
wire iffcq00txphaseshift180done;
wire iffcq00phyesmadaptationsave;
wire iffcq00rxdelayalignprogress;
wire iffcq00txdelayalignprogress;
wire iffcq00rxphasedelayresetdone;
wire iffcq00txphasedelayresetdone;
wire iffcq00txethernetstattxlocalfault;

wire [7:0]  iffcq00rxrate;
wire [7:0]  iffcq00txrate;
wire[127:0] iffcq00rxdata;
wire[127:0] iffcq00txdata;
wire [15:0] iffcq00rxctrl0;
wire [15:0] iffcq00rxctrl1;
wire [15:0] iffcq00txctrl0;
wire [15:0] iffcq00txctrl1;
wire [31:0] iffcq00dmonout;
wire [7:0]  iffcq00rxctrl2;
wire [7:0]  iffcq00rxctrl3;
wire [7:0]  iffcq00txctrl2;
wire [1:0]  iffcq00txdeemph;
wire [11:0] iffcq00bufgtdiv;
wire [15:0] iffcq00pinrsrvd;
wire [2:0]  iffcq00loopback;
wire [2:0]  iffcq00rxstatus;
wire [2:0]  iffcq00txmargin;
wire [4:0]  iffcq00txdrvamp;
wire [4:0]  iffcq00txemppos;
wire [4:0]  iffcq00txemppre;
wire [5:0]  iffcq00rxheader;
wire [5:0]  iffcq00txheader;
wire [1:0]  iffcq00refclkpma;
wire [15:0] iffcq00pcsrsvdin;
wire [3:0]  iffcq00rxprbssel;
wire [3:0]  iffcq00txprbssel;
wire [4:0]  iffcq00rxchbondi;
wire [4:0]  iffcq00rxchbondo;
wire [6:0]  iffcq00txempmain;
wire [1:0]  iffcq00rxckcorcnt;
wire [15:0] iffcq00pcsrsvdout;
wire [15:0] iffcq00pinrsrvdas;
wire [6:0]  iffcq00txsequence;
wire [1:0]  iffcq00rxdatavalid;
wire [1:0]  iffcq00rxpowerdown;
wire [1:0]  iffcq00rxresetmode;
wire [1:0]  iffcq00txbufstatus;
wire [1:0]  iffcq00txpowerdown;
wire [1:0]  iffcq00txresetmode;
wire [2:0]  iffcq00rxbufstatus;
wire [3:0]  iffcq00bufgtcemask;
wire [4:0]  iffcq00stepsizeppm;
wire [1:0]  iffcq00rxstartofseq;
wire [3:0]  iffcq00bufgtrstmask;
wire [1:0]  iffcq00rxheadervalid;
wire [2:0]  iffcq00txpmaresetmask;
wire [4:0]  iffcq00rxpcsresetmask;
wire [6:0]  iffcq00rxpmaresetmask;
wire [1:0]  iffcq00rxdapiresetmask;
wire [1:0]  iffcq00txdapiresetmask;
wire [1:0]  iffcq00rxchicoresetmask;
wire [1:0]  iffcq00txchicoresetmask;
wire [7:0]  iffcq00rxethernetstatout;

wire iffcq01enppm;
wire iffcq01perstb;
wire iffcq01bufgtce;
wire iffcq01cdrhold;
wire iffcq01cdrlock;
wire iffcq01dmonclk;
wire iffcq01rxlpmen;
wire iffcq01rxpkdet;
wire iffcq01rxqpien;
wire iffcq01rxslide;
wire iffcq01rxvalid;
wire iffcq01tstclk0;
wire iffcq01tstclk1;
wire iffcq01txswing;
wire iffcq01bufgtrst;
wire iffcq01cdrovren;
wire iffcq01cfokdone;
wire iffcq01iloreset;
wire iffcq01phyready;
wire iffcq01rxlatclk;
wire iffcq01rxusrclk;
wire iffcq01rxusrrdy;
wire iffcq01txcomsas;
wire iffcq01txlatclk;
wire iffcq01txusrclk;
wire iffcq01txusrrdy;
wire iffcq01bsrserial;
wire iffcq01cdrfreqos;
wire iffcq01cdrstepsq;
wire iffcq01cdrstepsx;
wire iffcq01comsasdet;
wire iffcq01gtrxreset;
wire iffcq01gttxreset;
wire iffcq01phystatus;
wire iffcq01rxprbserr;
wire iffcq01rxqpisenn;
wire iffcq01rxqpisenp;
wire iffcq01txcominit;
wire iffcq01txcomwake;
wire iffcq01txdccdone;
wire iffcq01txinhibit;
wire iffcq01txqpisenn;
wire iffcq01txqpisenp;
wire iffcq01aptexthold;
wire iffcq01cdrbmcdreq;
wire iffcq01cdrphreset;
wire iffcq01cdrstepdir;
wire iffcq01cominitdet;
wire iffcq01comwakedet;
wire iffcq01rxcommadet;
wire iffcq01rxelecidle;
wire iffcq01rxoobreset;
wire iffcq01rxpolarity;
wire iffcq01rxsliderdy;
wire iffcq01rxslipdone;
wire iffcq01rxsyncdone;
wire iffcq01txelecidle;
wire iffcq01txpolarity;
wire iffcq01txserpwrdn;
wire iffcq01txsyncdone;
wire iffcq01aptoverwren;
wire iffcq01cdrincpctrl;
wire iffcq01ckpinrsrvd0;
wire iffcq01ckpinrsrvd1;
wire iffcq01cssdstopclk;
wire iffcq01rxcdrphdone;
wire iffcq01rxdapireset;
wire iffcq01rxoutpcsclk;
wire iffcq01rxresetdone;
wire iffcq01rxsyncallin;
wire iffcq01txcomfinish;
wire iffcq01txdapireset;
wire iffcq01txoneszeros;
wire iffcq01txoutpcsclk;
wire iffcq01txqpibiasen;
wire iffcq01txqpiweakpu;
wire iffcq01txresetdone;
wire iffcq01txsyncallin;
wire iffcq01eyescanreset;
wire iffcq01hsdppcsreset;
wire iffcq01iloresetdone;
wire iffcq01iloresetmask;
wire iffcq01rxeqtraining;
wire iffcq01rxphdlyreset;
wire iffcq01rxprbslocked;
wire iffcq01txphdlyreset;
wire iffcq01dmonfiforeset;
wire iffcq01rxbyterealign;
wire iffcq01rxchanbondseq;
wire iffcq01rxchanrealign;
wire iffcq01rxchisaligned;
wire iffcq01rxgearboxslip;
wire iffcq01rxmldchainreq;
wire iffcq01rxtermination;
wire iffcq01txmldchainreq;
wire iffcq01txswingoutlow;
wire iffcq01eyescantrigger;
wire iffcq01resetexception;
wire iffcq01rxmldchaindone;
wire iffcq01rxphasealignpd;
wire iffcq01rxpmaresetdone;
wire iffcq01rxprbscntreset;
wire iffcq01rxprogdivreset;
wire iffcq01tcoclkfsmfrout;
wire iffcq01txchicooutrsvd;
wire iffcq01txmldchaindone;
wire iffcq01txpcsresetmask;
wire iffcq01txphasealignpd;
wire iffcq01txpmaresetdone;
wire iffcq01txprbsforceerr;
wire iffcq01txprogdivreset;
wire iffcq01txswingouthigh;
wire iffcq01rxbyteisaligned;
wire iffcq01rxdapicodereset;
wire iffcq01rxdapiresetdone;
wire iffcq01rxdelayalignerr;
wire iffcq01rxdelayalignreq;
wire iffcq01rxfinealigndone;
wire iffcq01rxphasealignerr;
wire iffcq01rxphasealignreq;
wire iffcq01txdapicodereset;
wire iffcq01txdapiresetdone;
wire iffcq01txdelayalignerr;
wire iffcq01txdelayalignreq;
wire iffcq01txphasealignerr;
wire iffcq01txphasealignreq;
wire iffcq01txtxpicodereset;
wire iffcq01eyescandataerror;
wire iffcq01rxdapicodeovrden;
wire iffcq01rxmlfinealignreq;
wire iffcq01rxphasealigndone;
wire iffcq01txdapicodeovrden;
wire iffcq01txphasealigndone;
wire iffcq01txtxpicodeovrden;
wire iffcq01xpipe5pipelineen;
wire iffcq01rxphasesetinitreq;
wire iffcq01txpausedelayalign;
wire iffcq01txphasesetinitreq;
wire iffcq01rxphasesetinitdone;
wire iffcq01rxphaseshift180req;
wire iffcq01rxprogdivresetdone;
wire iffcq01rxsimplexphystatus;
wire iffcq01txdetectrxloopback;
wire iffcq01txphasesetinitdone;
wire iffcq01txphaseshift180req;
wire iffcq01txprogdivresetdone;
wire iffcq01txsimplexphystatus;
wire iffcq01rxphaseshift180done;
wire iffcq01txphaseshift180done;
wire iffcq01phyesmadaptationsave;
wire iffcq01rxdelayalignprogress;
wire iffcq01txdelayalignprogress;
wire iffcq01rxphasedelayresetdone;
wire iffcq01txphasedelayresetdone;
wire iffcq01txethernetstattxlocalfault;

wire [7:0]  iffcq01rxrate;
wire [7:0]  iffcq01txrate;
wire[127:0] iffcq01rxdata;
wire[127:0] iffcq01txdata;
wire [15:0] iffcq01rxctrl0;
wire [15:0] iffcq01rxctrl1;
wire [15:0] iffcq01txctrl0;
wire [15:0] iffcq01txctrl1;
wire [31:0] iffcq01dmonout;
wire [7:0]  iffcq01rxctrl2;
wire [7:0]  iffcq01rxctrl3;
wire [7:0]  iffcq01txctrl2;
wire [1:0]  iffcq01txdeemph;
wire [11:0] iffcq01bufgtdiv;
wire [15:0] iffcq01pinrsrvd;
wire [2:0]  iffcq01loopback;
wire [2:0]  iffcq01rxstatus;
wire [2:0]  iffcq01txmargin;
wire [4:0]  iffcq01txdrvamp;
wire [4:0]  iffcq01txemppos;
wire [4:0]  iffcq01txemppre;
wire [5:0]  iffcq01rxheader;
wire [5:0]  iffcq01txheader;
wire [1:0]  iffcq01refclkpma;
wire [15:0] iffcq01pcsrsvdin;
wire [3:0]  iffcq01rxprbssel;
wire [3:0]  iffcq01txprbssel;
wire [4:0]  iffcq01rxchbondi;
wire [4:0]  iffcq01rxchbondo;
wire [6:0]  iffcq01txempmain;
wire [1:0]  iffcq01rxckcorcnt;
wire [15:0] iffcq01pcsrsvdout;
wire [15:0] iffcq01pinrsrvdas;
wire [6:0]  iffcq01txsequence;
wire [1:0]  iffcq01rxdatavalid;
wire [1:0]  iffcq01rxpowerdown;
wire [1:0]  iffcq01rxresetmode;
wire [1:0]  iffcq01txbufstatus;
wire [1:0]  iffcq01txpowerdown;
wire [1:0]  iffcq01txresetmode;
wire [2:0]  iffcq01rxbufstatus;
wire [3:0]  iffcq01bufgtcemask;
wire [4:0]  iffcq01stepsizeppm;
wire [1:0]  iffcq01rxstartofseq;
wire [3:0]  iffcq01bufgtrstmask;
wire [1:0]  iffcq01rxheadervalid;
wire [2:0]  iffcq01txpmaresetmask;
wire [4:0]  iffcq01rxpcsresetmask;
wire [6:0]  iffcq01rxpmaresetmask;
wire [1:0]  iffcq01rxdapiresetmask;
wire [1:0]  iffcq01txdapiresetmask;
wire [1:0]  iffcq01rxchicoresetmask;
wire [1:0]  iffcq01txchicoresetmask;
wire [7:0]  iffcq01rxethernetstatout;

wire iffcq02enppm;
wire iffcq02perstb;
wire iffcq02bufgtce;
wire iffcq02cdrhold;
wire iffcq02cdrlock;
wire iffcq02dmonclk;
wire iffcq02rxlpmen;
wire iffcq02rxpkdet;
wire iffcq02rxqpien;
wire iffcq02rxslide;
wire iffcq02rxvalid;
wire iffcq02tstclk0;
wire iffcq02tstclk1;
wire iffcq02txswing;
wire iffcq02bufgtrst;
wire iffcq02cdrovren;
wire iffcq02cfokdone;
wire iffcq02iloreset;
wire iffcq02phyready;
wire iffcq02rxlatclk;
wire iffcq02rxusrclk;
wire iffcq02rxusrrdy;
wire iffcq02txcomsas;
wire iffcq02txlatclk;
wire iffcq02txusrclk;
wire iffcq02txusrrdy;
wire iffcq02bsrserial;
wire iffcq02cdrfreqos;
wire iffcq02cdrstepsq;
wire iffcq02cdrstepsx;
wire iffcq02comsasdet;
wire iffcq02gtrxreset;
wire iffcq02gttxreset;
wire iffcq02phystatus;
wire iffcq02rxprbserr;
wire iffcq02rxqpisenn;
wire iffcq02rxqpisenp;
wire iffcq02txcominit;
wire iffcq02txcomwake;
wire iffcq02txdccdone;
wire iffcq02txinhibit;
wire iffcq02txqpisenn;
wire iffcq02txqpisenp;
wire iffcq02aptexthold;
wire iffcq02cdrbmcdreq;
wire iffcq02cdrphreset;
wire iffcq02cdrstepdir;
wire iffcq02cominitdet;
wire iffcq02comwakedet;
wire iffcq02rxcommadet;
wire iffcq02rxelecidle;
wire iffcq02rxoobreset;
wire iffcq02rxpolarity;
wire iffcq02rxsliderdy;
wire iffcq02rxslipdone;
wire iffcq02rxsyncdone;
wire iffcq02txelecidle;
wire iffcq02txpolarity;
wire iffcq02txserpwrdn;
wire iffcq02txsyncdone;
wire iffcq02aptoverwren;
wire iffcq02cdrincpctrl;
wire iffcq02ckpinrsrvd0;
wire iffcq02ckpinrsrvd1;
wire iffcq02cssdstopclk;
wire iffcq02rxcdrphdone;
wire iffcq02rxdapireset;
wire iffcq02rxoutpcsclk;
wire iffcq02rxresetdone;
wire iffcq02rxsyncallin;
wire iffcq02txcomfinish;
wire iffcq02txdapireset;
wire iffcq02txoneszeros;
wire iffcq02txoutpcsclk;
wire iffcq02txqpibiasen;
wire iffcq02txqpiweakpu;
wire iffcq02txresetdone;
wire iffcq02txsyncallin;
wire iffcq02eyescanreset;
wire iffcq02hsdppcsreset;
wire iffcq02iloresetdone;
wire iffcq02iloresetmask;
wire iffcq02rxeqtraining;
wire iffcq02rxphdlyreset;
wire iffcq02rxprbslocked;
wire iffcq02txphdlyreset;
wire iffcq02dmonfiforeset;
wire iffcq02rxbyterealign;
wire iffcq02rxchanbondseq;
wire iffcq02rxchanrealign;
wire iffcq02rxchisaligned;
wire iffcq02rxgearboxslip;
wire iffcq02rxmldchainreq;
wire iffcq02rxtermination;
wire iffcq02txmldchainreq;
wire iffcq02txswingoutlow;
wire iffcq02eyescantrigger;
wire iffcq02resetexception;
wire iffcq02rxmldchaindone;
wire iffcq02rxphasealignpd;
wire iffcq02rxpmaresetdone;
wire iffcq02rxprbscntreset;
wire iffcq02rxprogdivreset;
wire iffcq02tcoclkfsmfrout;
wire iffcq02txchicooutrsvd;
wire iffcq02txmldchaindone;
wire iffcq02txpcsresetmask;
wire iffcq02txphasealignpd;
wire iffcq02txpmaresetdone;
wire iffcq02txprbsforceerr;
wire iffcq02txprogdivreset;
wire iffcq02txswingouthigh;
wire iffcq02rxbyteisaligned;
wire iffcq02rxdapicodereset;
wire iffcq02rxdapiresetdone;
wire iffcq02rxdelayalignerr;
wire iffcq02rxdelayalignreq;
wire iffcq02rxfinealigndone;
wire iffcq02rxphasealignerr;
wire iffcq02rxphasealignreq;
wire iffcq02txdapicodereset;
wire iffcq02txdapiresetdone;
wire iffcq02txdelayalignerr;
wire iffcq02txdelayalignreq;
wire iffcq02txphasealignerr;
wire iffcq02txphasealignreq;
wire iffcq02txtxpicodereset;
wire iffcq02eyescandataerror;
wire iffcq02rxdapicodeovrden;
wire iffcq02rxmlfinealignreq;
wire iffcq02rxphasealigndone;
wire iffcq02txdapicodeovrden;
wire iffcq02txphasealigndone;
wire iffcq02txtxpicodeovrden;
wire iffcq02xpipe5pipelineen;
wire iffcq02rxphasesetinitreq;
wire iffcq02txpausedelayalign;
wire iffcq02txphasesetinitreq;
wire iffcq02rxphasesetinitdone;
wire iffcq02rxphaseshift180req;
wire iffcq02rxprogdivresetdone;
wire iffcq02rxsimplexphystatus;
wire iffcq02txdetectrxloopback;
wire iffcq02txphasesetinitdone;
wire iffcq02txphaseshift180req;
wire iffcq02txprogdivresetdone;
wire iffcq02txsimplexphystatus;
wire iffcq02rxphaseshift180done;
wire iffcq02txphaseshift180done;
wire iffcq02phyesmadaptationsave;
wire iffcq02rxdelayalignprogress;
wire iffcq02txdelayalignprogress;
wire iffcq02rxphasedelayresetdone;
wire iffcq02txphasedelayresetdone;
wire iffcq02txethernetstattxlocalfault;

wire [7:0]  iffcq02rxrate;
wire [7:0]  iffcq02txrate;
wire[127:0] iffcq02rxdata;
wire[127:0] iffcq02txdata;
wire [15:0] iffcq02rxctrl0;
wire [15:0] iffcq02rxctrl1;
wire [15:0] iffcq02txctrl0;
wire [15:0] iffcq02txctrl1;
wire [31:0] iffcq02dmonout;
wire [7:0]  iffcq02rxctrl2;
wire [7:0]  iffcq02rxctrl3;
wire [7:0]  iffcq02txctrl2;
wire [1:0]  iffcq02txdeemph;
wire [11:0] iffcq02bufgtdiv;
wire [15:0] iffcq02pinrsrvd;
wire [2:0]  iffcq02loopback;
wire [2:0]  iffcq02rxstatus;
wire [2:0]  iffcq02txmargin;
wire [4:0]  iffcq02txdrvamp;
wire [4:0]  iffcq02txemppos;
wire [4:0]  iffcq02txemppre;
wire [5:0]  iffcq02rxheader;
wire [5:0]  iffcq02txheader;
wire [1:0]  iffcq02refclkpma;
wire [15:0] iffcq02pcsrsvdin;
wire [3:0]  iffcq02rxprbssel;
wire [3:0]  iffcq02txprbssel;
wire [4:0]  iffcq02rxchbondi;
wire [4:0]  iffcq02rxchbondo;
wire [6:0]  iffcq02txempmain;
wire [1:0]  iffcq02rxckcorcnt;
wire [15:0] iffcq02pcsrsvdout;
wire [15:0] iffcq02pinrsrvdas;
wire [6:0]  iffcq02txsequence;
wire [1:0]  iffcq02rxdatavalid;
wire [1:0]  iffcq02rxpowerdown;
wire [1:0]  iffcq02rxresetmode;
wire [1:0]  iffcq02txbufstatus;
wire [1:0]  iffcq02txpowerdown;
wire [1:0]  iffcq02txresetmode;
wire [2:0]  iffcq02rxbufstatus;
wire [3:0]  iffcq02bufgtcemask;
wire [4:0]  iffcq02stepsizeppm;
wire [1:0]  iffcq02rxstartofseq;
wire [3:0]  iffcq02bufgtrstmask;
wire [1:0]  iffcq02rxheadervalid;
wire [2:0]  iffcq02txpmaresetmask;
wire [4:0]  iffcq02rxpcsresetmask;
wire [6:0]  iffcq02rxpmaresetmask;
wire [1:0]  iffcq02rxdapiresetmask;
wire [1:0]  iffcq02txdapiresetmask;
wire [1:0]  iffcq02rxchicoresetmask;
wire [1:0]  iffcq02txchicoresetmask;
wire [7:0]  iffcq02rxethernetstatout;

wire iffcq03enppm;
wire iffcq03perstb;
wire iffcq03bufgtce;
wire iffcq03cdrhold;
wire iffcq03cdrlock;
wire iffcq03dmonclk;
wire iffcq03rxlpmen;
wire iffcq03rxpkdet;
wire iffcq03rxqpien;
wire iffcq03rxslide;
wire iffcq03rxvalid;
wire iffcq03tstclk0;
wire iffcq03tstclk1;
wire iffcq03txswing;
wire iffcq03bufgtrst;
wire iffcq03cdrovren;
wire iffcq03cfokdone;
wire iffcq03iloreset;
wire iffcq03phyready;
wire iffcq03rxlatclk;
wire iffcq03rxusrclk;
wire iffcq03rxusrrdy;
wire iffcq03txcomsas;
wire iffcq03txlatclk;
wire iffcq03txusrclk;
wire iffcq03txusrrdy;
wire iffcq03bsrserial;
wire iffcq03cdrfreqos;
wire iffcq03cdrstepsq;
wire iffcq03cdrstepsx;
wire iffcq03comsasdet;
wire iffcq03gtrxreset;
wire iffcq03gttxreset;
wire iffcq03phystatus;
wire iffcq03rxprbserr;
wire iffcq03rxqpisenn;
wire iffcq03rxqpisenp;
wire iffcq03txcominit;
wire iffcq03txcomwake;
wire iffcq03txdccdone;
wire iffcq03txinhibit;
wire iffcq03txqpisenn;
wire iffcq03txqpisenp;
wire iffcq03aptexthold;
wire iffcq03cdrbmcdreq;
wire iffcq03cdrphreset;
wire iffcq03cdrstepdir;
wire iffcq03cominitdet;
wire iffcq03comwakedet;
wire iffcq03rxcommadet;
wire iffcq03rxelecidle;
wire iffcq03rxoobreset;
wire iffcq03rxpolarity;
wire iffcq03rxsliderdy;
wire iffcq03rxslipdone;
wire iffcq03rxsyncdone;
wire iffcq03txelecidle;
wire iffcq03txpolarity;
wire iffcq03txserpwrdn;
wire iffcq03txsyncdone;
wire iffcq03aptoverwren;
wire iffcq03cdrincpctrl;
wire iffcq03ckpinrsrvd0;
wire iffcq03ckpinrsrvd1;
wire iffcq03cssdstopclk;
wire iffcq03rxcdrphdone;
wire iffcq03rxdapireset;
wire iffcq03rxoutpcsclk;
wire iffcq03rxresetdone;
wire iffcq03rxsyncallin;
wire iffcq03txcomfinish;
wire iffcq03txdapireset;
wire iffcq03txoneszeros;
wire iffcq03txoutpcsclk;
wire iffcq03txqpibiasen;
wire iffcq03txqpiweakpu;
wire iffcq03txresetdone;
wire iffcq03txsyncallin;
wire iffcq03eyescanreset;
wire iffcq03hsdppcsreset;
wire iffcq03iloresetdone;
wire iffcq03iloresetmask;
wire iffcq03rxeqtraining;
wire iffcq03rxphdlyreset;
wire iffcq03rxprbslocked;
wire iffcq03txphdlyreset;
wire iffcq03dmonfiforeset;
wire iffcq03rxbyterealign;
wire iffcq03rxchanbondseq;
wire iffcq03rxchanrealign;
wire iffcq03rxchisaligned;
wire iffcq03rxgearboxslip;
wire iffcq03rxmldchainreq;
wire iffcq03rxtermination;
wire iffcq03txmldchainreq;
wire iffcq03txswingoutlow;
wire iffcq03eyescantrigger;
wire iffcq03resetexception;
wire iffcq03rxmldchaindone;
wire iffcq03rxphasealignpd;
wire iffcq03rxpmaresetdone;
wire iffcq03rxprbscntreset;
wire iffcq03rxprogdivreset;
wire iffcq03tcoclkfsmfrout;
wire iffcq03txchicooutrsvd;
wire iffcq03txmldchaindone;
wire iffcq03txpcsresetmask;
wire iffcq03txphasealignpd;
wire iffcq03txpmaresetdone;
wire iffcq03txprbsforceerr;
wire iffcq03txprogdivreset;
wire iffcq03txswingouthigh;
wire iffcq03rxbyteisaligned;
wire iffcq03rxdapicodereset;
wire iffcq03rxdapiresetdone;
wire iffcq03rxdelayalignerr;
wire iffcq03rxdelayalignreq;
wire iffcq03rxfinealigndone;
wire iffcq03rxphasealignerr;
wire iffcq03rxphasealignreq;
wire iffcq03txdapicodereset;
wire iffcq03txdapiresetdone;
wire iffcq03txdelayalignerr;
wire iffcq03txdelayalignreq;
wire iffcq03txphasealignerr;
wire iffcq03txphasealignreq;
wire iffcq03txtxpicodereset;
wire iffcq03eyescandataerror;
wire iffcq03rxdapicodeovrden;
wire iffcq03rxmlfinealignreq;
wire iffcq03rxphasealigndone;
wire iffcq03txdapicodeovrden;
wire iffcq03txphasealigndone;
wire iffcq03txtxpicodeovrden;
wire iffcq03xpipe5pipelineen;
wire iffcq03rxphasesetinitreq;
wire iffcq03txpausedelayalign;
wire iffcq03txphasesetinitreq;
wire iffcq03rxphasesetinitdone;
wire iffcq03rxphaseshift180req;
wire iffcq03rxprogdivresetdone;
wire iffcq03rxsimplexphystatus;
wire iffcq03txdetectrxloopback;
wire iffcq03txphasesetinitdone;
wire iffcq03txphaseshift180req;
wire iffcq03txprogdivresetdone;
wire iffcq03txsimplexphystatus;
wire iffcq03rxphaseshift180done;
wire iffcq03txphaseshift180done;
wire iffcq03phyesmadaptationsave;
wire iffcq03rxdelayalignprogress;
wire iffcq03txdelayalignprogress;
wire iffcq03rxphasedelayresetdone;
wire iffcq03txphasedelayresetdone;
wire iffcq03txethernetstattxlocalfault;

wire [7:0]  iffcq03rxrate;
wire [7:0]  iffcq03txrate;
wire[127:0] iffcq03rxdata;
wire[127:0] iffcq03txdata;
wire [15:0] iffcq03rxctrl0;
wire [15:0] iffcq03rxctrl1;
wire [15:0] iffcq03txctrl0;
wire [15:0] iffcq03txctrl1;
wire [31:0] iffcq03dmonout;
wire [7:0]  iffcq03rxctrl2;
wire [7:0]  iffcq03rxctrl3;
wire [7:0]  iffcq03txctrl2;
wire [1:0]  iffcq03txdeemph;
wire [11:0] iffcq03bufgtdiv;
wire [15:0] iffcq03pinrsrvd;
wire [2:0]  iffcq03loopback;
wire [2:0]  iffcq03rxstatus;
wire [2:0]  iffcq03txmargin;
wire [4:0]  iffcq03txdrvamp;
wire [4:0]  iffcq03txemppos;
wire [4:0]  iffcq03txemppre;
wire [5:0]  iffcq03rxheader;
wire [5:0]  iffcq03txheader;
wire [1:0]  iffcq03refclkpma;
wire [15:0] iffcq03pcsrsvdin;
wire [3:0]  iffcq03rxprbssel;
wire [3:0]  iffcq03txprbssel;
wire [4:0]  iffcq03rxchbondi;
wire [4:0]  iffcq03rxchbondo;
wire [6:0]  iffcq03txempmain;
wire [1:0]  iffcq03rxckcorcnt;
wire [15:0] iffcq03pcsrsvdout;
wire [15:0] iffcq03pinrsrvdas;
wire [6:0]  iffcq03txsequence;
wire [1:0]  iffcq03rxdatavalid;
wire [1:0]  iffcq03rxpowerdown;
wire [1:0]  iffcq03rxresetmode;
wire [1:0]  iffcq03txbufstatus;
wire [1:0]  iffcq03txpowerdown;
wire [1:0]  iffcq03txresetmode;
wire [2:0]  iffcq03rxbufstatus;
wire [3:0]  iffcq03bufgtcemask;
wire [4:0]  iffcq03stepsizeppm;
wire [1:0]  iffcq03rxstartofseq;
wire [3:0]  iffcq03bufgtrstmask;
wire [1:0]  iffcq03rxheadervalid;
wire [2:0]  iffcq03txpmaresetmask;
wire [4:0]  iffcq03rxpcsresetmask;
wire [6:0]  iffcq03rxpmaresetmask;
wire [1:0]  iffcq03rxdapiresetmask;
wire [1:0]  iffcq03txdapiresetmask;
wire [1:0]  iffcq03rxchicoresetmask;
wire [1:0]  iffcq03txchicoresetmask;
wire [7:0]  iffcq03rxethernetstatout;

wire iffcq10enppm;
wire iffcq10perstb;
wire iffcq10bufgtce;
wire iffcq10cdrhold;
wire iffcq10cdrlock;
wire iffcq10dmonclk;
wire iffcq10rxlpmen;
wire iffcq10rxpkdet;
wire iffcq10rxqpien;
wire iffcq10rxslide;
wire iffcq10rxvalid;
wire iffcq10tstclk0;
wire iffcq10tstclk1;
wire iffcq10txswing;
wire iffcq10bufgtrst;
wire iffcq10cdrovren;
wire iffcq10cfokdone;
wire iffcq10iloreset;
wire iffcq10phyready;
wire iffcq10rxlatclk;
wire iffcq10rxusrclk;
wire iffcq10rxusrrdy;
wire iffcq10txcomsas;
wire iffcq10txlatclk;
wire iffcq10txusrclk;
wire iffcq10txusrrdy;
wire iffcq10bsrserial;
wire iffcq10cdrfreqos;
wire iffcq10cdrstepsq;
wire iffcq10cdrstepsx;
wire iffcq10comsasdet;
wire iffcq10gtrxreset;
wire iffcq10gttxreset;
wire iffcq10phystatus;
wire iffcq10rxprbserr;
wire iffcq10rxqpisenn;
wire iffcq10rxqpisenp;
wire iffcq10txcominit;
wire iffcq10txcomwake;
wire iffcq10txdccdone;
wire iffcq10txinhibit;
wire iffcq10txqpisenn;
wire iffcq10txqpisenp;
wire iffcq10aptexthold;
wire iffcq10cdrbmcdreq;
wire iffcq10cdrphreset;
wire iffcq10cdrstepdir;
wire iffcq10cominitdet;
wire iffcq10comwakedet;
wire iffcq10rxcommadet;
wire iffcq10rxelecidle;
wire iffcq10rxoobreset;
wire iffcq10rxpolarity;
wire iffcq10rxsliderdy;
wire iffcq10rxslipdone;
wire iffcq10rxsyncdone;
wire iffcq10txelecidle;
wire iffcq10txpolarity;
wire iffcq10txserpwrdn;
wire iffcq10txsyncdone;
wire iffcq10aptoverwren;
wire iffcq10cdrincpctrl;
wire iffcq10ckpinrsrvd0;
wire iffcq10ckpinrsrvd1;
wire iffcq10cssdstopclk;
wire iffcq10rxcdrphdone;
wire iffcq10rxdapireset;
wire iffcq10rxoutpcsclk;
wire iffcq10rxresetdone;
wire iffcq10rxsyncallin;
wire iffcq10txcomfinish;
wire iffcq10txdapireset;
wire iffcq10txoneszeros;
wire iffcq10txoutpcsclk;
wire iffcq10txqpibiasen;
wire iffcq10txqpiweakpu;
wire iffcq10txresetdone;
wire iffcq10txsyncallin;
wire iffcq10eyescanreset;
wire iffcq10hsdppcsreset;
wire iffcq10iloresetdone;
wire iffcq10iloresetmask;
wire iffcq10rxeqtraining;
wire iffcq10rxphdlyreset;
wire iffcq10rxprbslocked;
wire iffcq10txphdlyreset;
wire iffcq10dmonfiforeset;
wire iffcq10rxbyterealign;
wire iffcq10rxchanbondseq;
wire iffcq10rxchanrealign;
wire iffcq10rxchisaligned;
wire iffcq10rxgearboxslip;
wire iffcq10rxmldchainreq;
wire iffcq10rxtermination;
wire iffcq10txmldchainreq;
wire iffcq10txswingoutlow;
wire iffcq10eyescantrigger;
wire iffcq10resetexception;
wire iffcq10rxmldchaindone;
wire iffcq10rxphasealignpd;
wire iffcq10rxpmaresetdone;
wire iffcq10rxprbscntreset;
wire iffcq10rxprogdivreset;
wire iffcq10tcoclkfsmfrout;
wire iffcq10txchicooutrsvd;
wire iffcq10txmldchaindone;
wire iffcq10txpcsresetmask;
wire iffcq10txphasealignpd;
wire iffcq10txpmaresetdone;
wire iffcq10txprbsforceerr;
wire iffcq10txprogdivreset;
wire iffcq10txswingouthigh;
wire iffcq10rxbyteisaligned;
wire iffcq10rxdapicodereset;
wire iffcq10rxdapiresetdone;
wire iffcq10rxdelayalignerr;
wire iffcq10rxdelayalignreq;
wire iffcq10rxfinealigndone;
wire iffcq10rxphasealignerr;
wire iffcq10rxphasealignreq;
wire iffcq10txdapicodereset;
wire iffcq10txdapiresetdone;
wire iffcq10txdelayalignerr;
wire iffcq10txdelayalignreq;
wire iffcq10txphasealignerr;
wire iffcq10txphasealignreq;
wire iffcq10txtxpicodereset;
wire iffcq10eyescandataerror;
wire iffcq10rxdapicodeovrden;
wire iffcq10rxmlfinealignreq;
wire iffcq10rxphasealigndone;
wire iffcq10txdapicodeovrden;
wire iffcq10txphasealigndone;
wire iffcq10txtxpicodeovrden;
wire iffcq10xpipe5pipelineen;
wire iffcq10rxphasesetinitreq;
wire iffcq10txpausedelayalign;
wire iffcq10txphasesetinitreq;
wire iffcq10rxphasesetinitdone;
wire iffcq10rxphaseshift180req;
wire iffcq10rxprogdivresetdone;
wire iffcq10rxsimplexphystatus;
wire iffcq10txdetectrxloopback;
wire iffcq10txphasesetinitdone;
wire iffcq10txphaseshift180req;
wire iffcq10txprogdivresetdone;
wire iffcq10txsimplexphystatus;
wire iffcq10rxphaseshift180done;
wire iffcq10txphaseshift180done;
wire iffcq10phyesmadaptationsave;
wire iffcq10rxdelayalignprogress;
wire iffcq10txdelayalignprogress;
wire iffcq10rxphasedelayresetdone;
wire iffcq10txphasedelayresetdone;
wire iffcq10txethernetstattxlocalfault;

wire [7:0]  iffcq10rxrate;
wire [7:0]  iffcq10txrate;
wire[127:0] iffcq10rxdata;
wire[127:0] iffcq10txdata;
wire [15:0] iffcq10rxctrl0;
wire [15:0] iffcq10rxctrl1;
wire [15:0] iffcq10txctrl0;
wire [15:0] iffcq10txctrl1;
wire [31:0] iffcq10dmonout;
wire [7:0]  iffcq10rxctrl2;
wire [7:0]  iffcq10rxctrl3;
wire [7:0]  iffcq10txctrl2;
wire [1:0]  iffcq10txdeemph;
wire [11:0] iffcq10bufgtdiv;
wire [15:0] iffcq10pinrsrvd;
wire [2:0]  iffcq10loopback;
wire [2:0]  iffcq10rxstatus;
wire [2:0]  iffcq10txmargin;
wire [4:0]  iffcq10txdrvamp;
wire [4:0]  iffcq10txemppos;
wire [4:0]  iffcq10txemppre;
wire [5:0]  iffcq10rxheader;
wire [5:0]  iffcq10txheader;
wire [1:0]  iffcq10refclkpma;
wire [15:0] iffcq10pcsrsvdin;
wire [3:0]  iffcq10rxprbssel;
wire [3:0]  iffcq10txprbssel;
wire [4:0]  iffcq10rxchbondi;
wire [4:0]  iffcq10rxchbondo;
wire [6:0]  iffcq10txempmain;
wire [1:0]  iffcq10rxckcorcnt;
wire [15:0] iffcq10pcsrsvdout;
wire [15:0] iffcq10pinrsrvdas;
wire [6:0]  iffcq10txsequence;
wire [1:0]  iffcq10rxdatavalid;
wire [1:0]  iffcq10rxpowerdown;
wire [1:0]  iffcq10rxresetmode;
wire [1:0]  iffcq10txbufstatus;
wire [1:0]  iffcq10txpowerdown;
wire [1:0]  iffcq10txresetmode;
wire [2:0]  iffcq10rxbufstatus;
wire [3:0]  iffcq10bufgtcemask;
wire [4:0]  iffcq10stepsizeppm;
wire [1:0]  iffcq10rxstartofseq;
wire [3:0]  iffcq10bufgtrstmask;
wire [1:0]  iffcq10rxheadervalid;
wire [2:0]  iffcq10txpmaresetmask;
wire [4:0]  iffcq10rxpcsresetmask;
wire [6:0]  iffcq10rxpmaresetmask;
wire [1:0]  iffcq10rxdapiresetmask;
wire [1:0]  iffcq10txdapiresetmask;
wire [1:0]  iffcq10rxchicoresetmask;
wire [1:0]  iffcq10txchicoresetmask;
wire [7:0]  iffcq10rxethernetstatout;

wire iffcq11enppm;
wire iffcq11perstb;
wire iffcq11bufgtce;
wire iffcq11cdrhold;
wire iffcq11cdrlock;
wire iffcq11dmonclk;
wire iffcq11rxlpmen;
wire iffcq11rxpkdet;
wire iffcq11rxqpien;
wire iffcq11rxslide;
wire iffcq11rxvalid;
wire iffcq11tstclk0;
wire iffcq11tstclk1;
wire iffcq11txswing;
wire iffcq11bufgtrst;
wire iffcq11cdrovren;
wire iffcq11cfokdone;
wire iffcq11iloreset;
wire iffcq11phyready;
wire iffcq11rxlatclk;
wire iffcq11rxusrclk;
wire iffcq11rxusrrdy;
wire iffcq11txcomsas;
wire iffcq11txlatclk;
wire iffcq11txusrclk;
wire iffcq11txusrrdy;
wire iffcq11bsrserial;
wire iffcq11cdrfreqos;
wire iffcq11cdrstepsq;
wire iffcq11cdrstepsx;
wire iffcq11comsasdet;
wire iffcq11gtrxreset;
wire iffcq11gttxreset;
wire iffcq11phystatus;
wire iffcq11rxprbserr;
wire iffcq11rxqpisenn;
wire iffcq11rxqpisenp;
wire iffcq11txcominit;
wire iffcq11txcomwake;
wire iffcq11txdccdone;
wire iffcq11txinhibit;
wire iffcq11txqpisenn;
wire iffcq11txqpisenp;
wire iffcq11aptexthold;
wire iffcq11cdrbmcdreq;
wire iffcq11cdrphreset;
wire iffcq11cdrstepdir;
wire iffcq11cominitdet;
wire iffcq11comwakedet;
wire iffcq11rxcommadet;
wire iffcq11rxelecidle;
wire iffcq11rxoobreset;
wire iffcq11rxpolarity;
wire iffcq11rxsliderdy;
wire iffcq11rxslipdone;
wire iffcq11rxsyncdone;
wire iffcq11txelecidle;
wire iffcq11txpolarity;
wire iffcq11txserpwrdn;
wire iffcq11txsyncdone;
wire iffcq11aptoverwren;
wire iffcq11cdrincpctrl;
wire iffcq11ckpinrsrvd0;
wire iffcq11ckpinrsrvd1;
wire iffcq11cssdstopclk;
wire iffcq11rxcdrphdone;
wire iffcq11rxdapireset;
wire iffcq11rxoutpcsclk;
wire iffcq11rxresetdone;
wire iffcq11rxsyncallin;
wire iffcq11txcomfinish;
wire iffcq11txdapireset;
wire iffcq11txoneszeros;
wire iffcq11txoutpcsclk;
wire iffcq11txqpibiasen;
wire iffcq11txqpiweakpu;
wire iffcq11txresetdone;
wire iffcq11txsyncallin;
wire iffcq11eyescanreset;
wire iffcq11hsdppcsreset;
wire iffcq11iloresetdone;
wire iffcq11iloresetmask;
wire iffcq11rxeqtraining;
wire iffcq11rxphdlyreset;
wire iffcq11rxprbslocked;
wire iffcq11txphdlyreset;
wire iffcq11dmonfiforeset;
wire iffcq11rxbyterealign;
wire iffcq11rxchanbondseq;
wire iffcq11rxchanrealign;
wire iffcq11rxchisaligned;
wire iffcq11rxgearboxslip;
wire iffcq11rxmldchainreq;
wire iffcq11rxtermination;
wire iffcq11txmldchainreq;
wire iffcq11txswingoutlow;
wire iffcq11eyescantrigger;
wire iffcq11resetexception;
wire iffcq11rxmldchaindone;
wire iffcq11rxphasealignpd;
wire iffcq11rxpmaresetdone;
wire iffcq11rxprbscntreset;
wire iffcq11rxprogdivreset;
wire iffcq11tcoclkfsmfrout;
wire iffcq11txchicooutrsvd;
wire iffcq11txmldchaindone;
wire iffcq11txpcsresetmask;
wire iffcq11txphasealignpd;
wire iffcq11txpmaresetdone;
wire iffcq11txprbsforceerr;
wire iffcq11txprogdivreset;
wire iffcq11txswingouthigh;
wire iffcq11rxbyteisaligned;
wire iffcq11rxdapicodereset;
wire iffcq11rxdapiresetdone;
wire iffcq11rxdelayalignerr;
wire iffcq11rxdelayalignreq;
wire iffcq11rxfinealigndone;
wire iffcq11rxphasealignerr;
wire iffcq11rxphasealignreq;
wire iffcq11txdapicodereset;
wire iffcq11txdapiresetdone;
wire iffcq11txdelayalignerr;
wire iffcq11txdelayalignreq;
wire iffcq11txphasealignerr;
wire iffcq11txphasealignreq;
wire iffcq11txtxpicodereset;
wire iffcq11eyescandataerror;
wire iffcq11rxdapicodeovrden;
wire iffcq11rxmlfinealignreq;
wire iffcq11rxphasealigndone;
wire iffcq11txdapicodeovrden;
wire iffcq11txphasealigndone;
wire iffcq11txtxpicodeovrden;
wire iffcq11xpipe5pipelineen;
wire iffcq11rxphasesetinitreq;
wire iffcq11txpausedelayalign;
wire iffcq11txphasesetinitreq;
wire iffcq11rxphasesetinitdone;
wire iffcq11rxphaseshift180req;
wire iffcq11rxprogdivresetdone;
wire iffcq11rxsimplexphystatus;
wire iffcq11txdetectrxloopback;
wire iffcq11txphasesetinitdone;
wire iffcq11txphaseshift180req;
wire iffcq11txprogdivresetdone;
wire iffcq11txsimplexphystatus;
wire iffcq11rxphaseshift180done;
wire iffcq11txphaseshift180done;
wire iffcq11phyesmadaptationsave;
wire iffcq11rxdelayalignprogress;
wire iffcq11txdelayalignprogress;
wire iffcq11rxphasedelayresetdone;
wire iffcq11txphasedelayresetdone;
wire iffcq11txethernetstattxlocalfault;

wire [7:0]  iffcq11rxrate;
wire [7:0]  iffcq11txrate;
wire[127:0] iffcq11rxdata;
wire[127:0] iffcq11txdata;
wire [15:0] iffcq11rxctrl0;
wire [15:0] iffcq11rxctrl1;
wire [15:0] iffcq11txctrl0;
wire [15:0] iffcq11txctrl1;
wire [31:0] iffcq11dmonout;
wire [7:0]  iffcq11rxctrl2;
wire [7:0]  iffcq11rxctrl3;
wire [7:0]  iffcq11txctrl2;
wire [1:0]  iffcq11txdeemph;
wire [11:0] iffcq11bufgtdiv;
wire [15:0] iffcq11pinrsrvd;
wire [2:0]  iffcq11loopback;
wire [2:0]  iffcq11rxstatus;
wire [2:0]  iffcq11txmargin;
wire [4:0]  iffcq11txdrvamp;
wire [4:0]  iffcq11txemppos;
wire [4:0]  iffcq11txemppre;
wire [5:0]  iffcq11rxheader;
wire [5:0]  iffcq11txheader;
wire [1:0]  iffcq11refclkpma;
wire [15:0] iffcq11pcsrsvdin;
wire [3:0]  iffcq11rxprbssel;
wire [3:0]  iffcq11txprbssel;
wire [4:0]  iffcq11rxchbondi;
wire [4:0]  iffcq11rxchbondo;
wire [6:0]  iffcq11txempmain;
wire [1:0]  iffcq11rxckcorcnt;
wire [15:0] iffcq11pcsrsvdout;
wire [15:0] iffcq11pinrsrvdas;
wire [6:0]  iffcq11txsequence;
wire [1:0]  iffcq11rxdatavalid;
wire [1:0]  iffcq11rxpowerdown;
wire [1:0]  iffcq11rxresetmode;
wire [1:0]  iffcq11txbufstatus;
wire [1:0]  iffcq11txpowerdown;
wire [1:0]  iffcq11txresetmode;
wire [2:0]  iffcq11rxbufstatus;
wire [3:0]  iffcq11bufgtcemask;
wire [4:0]  iffcq11stepsizeppm;
wire [1:0]  iffcq11rxstartofseq;
wire [3:0]  iffcq11bufgtrstmask;
wire [1:0]  iffcq11rxheadervalid;
wire [2:0]  iffcq11txpmaresetmask;
wire [4:0]  iffcq11rxpcsresetmask;
wire [6:0]  iffcq11rxpmaresetmask;
wire [1:0]  iffcq11rxdapiresetmask;
wire [1:0]  iffcq11txdapiresetmask;
wire [1:0]  iffcq11rxchicoresetmask;
wire [1:0]  iffcq11txchicoresetmask;
wire [7:0]  iffcq11rxethernetstatout;

wire iffcq12enppm;
wire iffcq12perstb;
wire iffcq12bufgtce;
wire iffcq12cdrhold;
wire iffcq12cdrlock;
wire iffcq12dmonclk;
wire iffcq12rxlpmen;
wire iffcq12rxpkdet;
wire iffcq12rxqpien;
wire iffcq12rxslide;
wire iffcq12rxvalid;
wire iffcq12tstclk0;
wire iffcq12tstclk1;
wire iffcq12txswing;
wire iffcq12bufgtrst;
wire iffcq12cdrovren;
wire iffcq12cfokdone;
wire iffcq12iloreset;
wire iffcq12phyready;
wire iffcq12rxlatclk;
wire iffcq12rxusrclk;
wire iffcq12rxusrrdy;
wire iffcq12txcomsas;
wire iffcq12txlatclk;
wire iffcq12txusrclk;
wire iffcq12txusrrdy;
wire iffcq12bsrserial;
wire iffcq12cdrfreqos;
wire iffcq12cdrstepsq;
wire iffcq12cdrstepsx;
wire iffcq12comsasdet;
wire iffcq12gtrxreset;
wire iffcq12gttxreset;
wire iffcq12phystatus;
wire iffcq12rxprbserr;
wire iffcq12rxqpisenn;
wire iffcq12rxqpisenp;
wire iffcq12txcominit;
wire iffcq12txcomwake;
wire iffcq12txdccdone;
wire iffcq12txinhibit;
wire iffcq12txqpisenn;
wire iffcq12txqpisenp;
wire iffcq12aptexthold;
wire iffcq12cdrbmcdreq;
wire iffcq12cdrphreset;
wire iffcq12cdrstepdir;
wire iffcq12cominitdet;
wire iffcq12comwakedet;
wire iffcq12rxcommadet;
wire iffcq12rxelecidle;
wire iffcq12rxoobreset;
wire iffcq12rxpolarity;
wire iffcq12rxsliderdy;
wire iffcq12rxslipdone;
wire iffcq12rxsyncdone;
wire iffcq12txelecidle;
wire iffcq12txpolarity;
wire iffcq12txserpwrdn;
wire iffcq12txsyncdone;
wire iffcq12aptoverwren;
wire iffcq12cdrincpctrl;
wire iffcq12ckpinrsrvd0;
wire iffcq12ckpinrsrvd1;
wire iffcq12cssdstopclk;
wire iffcq12rxcdrphdone;
wire iffcq12rxdapireset;
wire iffcq12rxoutpcsclk;
wire iffcq12rxresetdone;
wire iffcq12rxsyncallin;
wire iffcq12txcomfinish;
wire iffcq12txdapireset;
wire iffcq12txoneszeros;
wire iffcq12txoutpcsclk;
wire iffcq12txqpibiasen;
wire iffcq12txqpiweakpu;
wire iffcq12txresetdone;
wire iffcq12txsyncallin;
wire iffcq12eyescanreset;
wire iffcq12hsdppcsreset;
wire iffcq12iloresetdone;
wire iffcq12iloresetmask;
wire iffcq12rxeqtraining;
wire iffcq12rxphdlyreset;
wire iffcq12rxprbslocked;
wire iffcq12txphdlyreset;
wire iffcq12dmonfiforeset;
wire iffcq12rxbyterealign;
wire iffcq12rxchanbondseq;
wire iffcq12rxchanrealign;
wire iffcq12rxchisaligned;
wire iffcq12rxgearboxslip;
wire iffcq12rxmldchainreq;
wire iffcq12rxtermination;
wire iffcq12txmldchainreq;
wire iffcq12txswingoutlow;
wire iffcq12eyescantrigger;
wire iffcq12resetexception;
wire iffcq12rxmldchaindone;
wire iffcq12rxphasealignpd;
wire iffcq12rxpmaresetdone;
wire iffcq12rxprbscntreset;
wire iffcq12rxprogdivreset;
wire iffcq12tcoclkfsmfrout;
wire iffcq12txchicooutrsvd;
wire iffcq12txmldchaindone;
wire iffcq12txpcsresetmask;
wire iffcq12txphasealignpd;
wire iffcq12txpmaresetdone;
wire iffcq12txprbsforceerr;
wire iffcq12txprogdivreset;
wire iffcq12txswingouthigh;
wire iffcq12rxbyteisaligned;
wire iffcq12rxdapicodereset;
wire iffcq12rxdapiresetdone;
wire iffcq12rxdelayalignerr;
wire iffcq12rxdelayalignreq;
wire iffcq12rxfinealigndone;
wire iffcq12rxphasealignerr;
wire iffcq12rxphasealignreq;
wire iffcq12txdapicodereset;
wire iffcq12txdapiresetdone;
wire iffcq12txdelayalignerr;
wire iffcq12txdelayalignreq;
wire iffcq12txphasealignerr;
wire iffcq12txphasealignreq;
wire iffcq12txtxpicodereset;
wire iffcq12eyescandataerror;
wire iffcq12rxdapicodeovrden;
wire iffcq12rxmlfinealignreq;
wire iffcq12rxphasealigndone;
wire iffcq12txdapicodeovrden;
wire iffcq12txphasealigndone;
wire iffcq12txtxpicodeovrden;
wire iffcq12xpipe5pipelineen;
wire iffcq12rxphasesetinitreq;
wire iffcq12txpausedelayalign;
wire iffcq12txphasesetinitreq;
wire iffcq12rxphasesetinitdone;
wire iffcq12rxphaseshift180req;
wire iffcq12rxprogdivresetdone;
wire iffcq12rxsimplexphystatus;
wire iffcq12txdetectrxloopback;
wire iffcq12txphasesetinitdone;
wire iffcq12txphaseshift180req;
wire iffcq12txprogdivresetdone;
wire iffcq12txsimplexphystatus;
wire iffcq12rxphaseshift180done;
wire iffcq12txphaseshift180done;
wire iffcq12phyesmadaptationsave;
wire iffcq12rxdelayalignprogress;
wire iffcq12txdelayalignprogress;
wire iffcq12rxphasedelayresetdone;
wire iffcq12txphasedelayresetdone;
wire iffcq12txethernetstattxlocalfault;

wire [7:0]  iffcq12rxrate;
wire [7:0]  iffcq12txrate;
wire[127:0] iffcq12rxdata;
wire[127:0] iffcq12txdata;
wire [15:0] iffcq12rxctrl0;
wire [15:0] iffcq12rxctrl1;
wire [15:0] iffcq12txctrl0;
wire [15:0] iffcq12txctrl1;
wire [31:0] iffcq12dmonout;
wire [7:0]  iffcq12rxctrl2;
wire [7:0]  iffcq12rxctrl3;
wire [7:0]  iffcq12txctrl2;
wire [1:0]  iffcq12txdeemph;
wire [11:0] iffcq12bufgtdiv;
wire [15:0] iffcq12pinrsrvd;
wire [2:0]  iffcq12loopback;
wire [2:0]  iffcq12rxstatus;
wire [2:0]  iffcq12txmargin;
wire [4:0]  iffcq12txdrvamp;
wire [4:0]  iffcq12txemppos;
wire [4:0]  iffcq12txemppre;
wire [5:0]  iffcq12rxheader;
wire [5:0]  iffcq12txheader;
wire [1:0]  iffcq12refclkpma;
wire [15:0] iffcq12pcsrsvdin;
wire [3:0]  iffcq12rxprbssel;
wire [3:0]  iffcq12txprbssel;
wire [4:0]  iffcq12rxchbondi;
wire [4:0]  iffcq12rxchbondo;
wire [6:0]  iffcq12txempmain;
wire [1:0]  iffcq12rxckcorcnt;
wire [15:0] iffcq12pcsrsvdout;
wire [15:0] iffcq12pinrsrvdas;
wire [6:0]  iffcq12txsequence;
wire [1:0]  iffcq12rxdatavalid;
wire [1:0]  iffcq12rxpowerdown;
wire [1:0]  iffcq12rxresetmode;
wire [1:0]  iffcq12txbufstatus;
wire [1:0]  iffcq12txpowerdown;
wire [1:0]  iffcq12txresetmode;
wire [2:0]  iffcq12rxbufstatus;
wire [3:0]  iffcq12bufgtcemask;
wire [4:0]  iffcq12stepsizeppm;
wire [1:0]  iffcq12rxstartofseq;
wire [3:0]  iffcq12bufgtrstmask;
wire [1:0]  iffcq12rxheadervalid;
wire [2:0]  iffcq12txpmaresetmask;
wire [4:0]  iffcq12rxpcsresetmask;
wire [6:0]  iffcq12rxpmaresetmask;
wire [1:0]  iffcq12rxdapiresetmask;
wire [1:0]  iffcq12txdapiresetmask;
wire [1:0]  iffcq12rxchicoresetmask;
wire [1:0]  iffcq12txchicoresetmask;
wire [7:0]  iffcq12rxethernetstatout;

wire iffcq13enppm;
wire iffcq13perstb;
wire iffcq13bufgtce;
wire iffcq13cdrhold;
wire iffcq13cdrlock;
wire iffcq13dmonclk;
wire iffcq13rxlpmen;
wire iffcq13rxpkdet;
wire iffcq13rxqpien;
wire iffcq13rxslide;
wire iffcq13rxvalid;
wire iffcq13tstclk0;
wire iffcq13tstclk1;
wire iffcq13txswing;
wire iffcq13bufgtrst;
wire iffcq13cdrovren;
wire iffcq13cfokdone;
wire iffcq13iloreset;
wire iffcq13phyready;
wire iffcq13rxlatclk;
wire iffcq13rxusrclk;
wire iffcq13rxusrrdy;
wire iffcq13txcomsas;
wire iffcq13txlatclk;
wire iffcq13txusrclk;
wire iffcq13txusrrdy;
wire iffcq13bsrserial;
wire iffcq13cdrfreqos;
wire iffcq13cdrstepsq;
wire iffcq13cdrstepsx;
wire iffcq13comsasdet;
wire iffcq13gtrxreset;
wire iffcq13gttxreset;
wire iffcq13phystatus;
wire iffcq13rxprbserr;
wire iffcq13rxqpisenn;
wire iffcq13rxqpisenp;
wire iffcq13txcominit;
wire iffcq13txcomwake;
wire iffcq13txdccdone;
wire iffcq13txinhibit;
wire iffcq13txqpisenn;
wire iffcq13txqpisenp;
wire iffcq13aptexthold;
wire iffcq13cdrbmcdreq;
wire iffcq13cdrphreset;
wire iffcq13cdrstepdir;
wire iffcq13cominitdet;
wire iffcq13comwakedet;
wire iffcq13rxcommadet;
wire iffcq13rxelecidle;
wire iffcq13rxoobreset;
wire iffcq13rxpolarity;
wire iffcq13rxsliderdy;
wire iffcq13rxslipdone;
wire iffcq13rxsyncdone;
wire iffcq13txelecidle;
wire iffcq13txpolarity;
wire iffcq13txserpwrdn;
wire iffcq13txsyncdone;
wire iffcq13aptoverwren;
wire iffcq13cdrincpctrl;
wire iffcq13ckpinrsrvd0;
wire iffcq13ckpinrsrvd1;
wire iffcq13cssdstopclk;
wire iffcq13rxcdrphdone;
wire iffcq13rxdapireset;
wire iffcq13rxoutpcsclk;
wire iffcq13rxresetdone;
wire iffcq13rxsyncallin;
wire iffcq13txcomfinish;
wire iffcq13txdapireset;
wire iffcq13txoneszeros;
wire iffcq13txoutpcsclk;
wire iffcq13txqpibiasen;
wire iffcq13txqpiweakpu;
wire iffcq13txresetdone;
wire iffcq13txsyncallin;
wire iffcq13eyescanreset;
wire iffcq13hsdppcsreset;
wire iffcq13iloresetdone;
wire iffcq13iloresetmask;
wire iffcq13rxeqtraining;
wire iffcq13rxphdlyreset;
wire iffcq13rxprbslocked;
wire iffcq13txphdlyreset;
wire iffcq13dmonfiforeset;
wire iffcq13rxbyterealign;
wire iffcq13rxchanbondseq;
wire iffcq13rxchanrealign;
wire iffcq13rxchisaligned;
wire iffcq13rxgearboxslip;
wire iffcq13rxmldchainreq;
wire iffcq13rxtermination;
wire iffcq13txmldchainreq;
wire iffcq13txswingoutlow;
wire iffcq13eyescantrigger;
wire iffcq13resetexception;
wire iffcq13rxmldchaindone;
wire iffcq13rxphasealignpd;
wire iffcq13rxpmaresetdone;
wire iffcq13rxprbscntreset;
wire iffcq13rxprogdivreset;
wire iffcq13tcoclkfsmfrout;
wire iffcq13txchicooutrsvd;
wire iffcq13txmldchaindone;
wire iffcq13txpcsresetmask;
wire iffcq13txphasealignpd;
wire iffcq13txpmaresetdone;
wire iffcq13txprbsforceerr;
wire iffcq13txprogdivreset;
wire iffcq13txswingouthigh;
wire iffcq13rxbyteisaligned;
wire iffcq13rxdapicodereset;
wire iffcq13rxdapiresetdone;
wire iffcq13rxdelayalignerr;
wire iffcq13rxdelayalignreq;
wire iffcq13rxfinealigndone;
wire iffcq13rxphasealignerr;
wire iffcq13rxphasealignreq;
wire iffcq13txdapicodereset;
wire iffcq13txdapiresetdone;
wire iffcq13txdelayalignerr;
wire iffcq13txdelayalignreq;
wire iffcq13txphasealignerr;
wire iffcq13txphasealignreq;
wire iffcq13txtxpicodereset;
wire iffcq13eyescandataerror;
wire iffcq13rxdapicodeovrden;
wire iffcq13rxmlfinealignreq;
wire iffcq13rxphasealigndone;
wire iffcq13txdapicodeovrden;
wire iffcq13txphasealigndone;
wire iffcq13txtxpicodeovrden;
wire iffcq13xpipe5pipelineen;
wire iffcq13rxphasesetinitreq;
wire iffcq13txpausedelayalign;
wire iffcq13txphasesetinitreq;
wire iffcq13rxphasesetinitdone;
wire iffcq13rxphaseshift180req;
wire iffcq13rxprogdivresetdone;
wire iffcq13rxsimplexphystatus;
wire iffcq13txdetectrxloopback;
wire iffcq13txphasesetinitdone;
wire iffcq13txphaseshift180req;
wire iffcq13txprogdivresetdone;
wire iffcq13txsimplexphystatus;
wire iffcq13rxphaseshift180done;
wire iffcq13txphaseshift180done;
wire iffcq13phyesmadaptationsave;
wire iffcq13rxdelayalignprogress;
wire iffcq13txdelayalignprogress;
wire iffcq13rxphasedelayresetdone;
wire iffcq13txphasedelayresetdone;
wire iffcq13txethernetstattxlocalfault;

wire [7:0]  iffcq13rxrate;
wire [7:0]  iffcq13txrate;
wire[127:0] iffcq13rxdata;
wire[127:0] iffcq13txdata;
wire [15:0] iffcq13rxctrl0;
wire [15:0] iffcq13rxctrl1;
wire [15:0] iffcq13txctrl0;
wire [15:0] iffcq13txctrl1;
wire [31:0] iffcq13dmonout;
wire [7:0]  iffcq13rxctrl2;
wire [7:0]  iffcq13rxctrl3;
wire [7:0]  iffcq13txctrl2;
wire [1:0]  iffcq13txdeemph;
wire [11:0] iffcq13bufgtdiv;
wire [15:0] iffcq13pinrsrvd;
wire [2:0]  iffcq13loopback;
wire [2:0]  iffcq13rxstatus;
wire [2:0]  iffcq13txmargin;
wire [4:0]  iffcq13txdrvamp;
wire [4:0]  iffcq13txemppos;
wire [4:0]  iffcq13txemppre;
wire [5:0]  iffcq13rxheader;
wire [5:0]  iffcq13txheader;
wire [1:0]  iffcq13refclkpma;
wire [15:0] iffcq13pcsrsvdin;
wire [3:0]  iffcq13rxprbssel;
wire [3:0]  iffcq13txprbssel;
wire [4:0]  iffcq13rxchbondi;
wire [4:0]  iffcq13rxchbondo;
wire [6:0]  iffcq13txempmain;
wire [1:0]  iffcq13rxckcorcnt;
wire [15:0] iffcq13pcsrsvdout;
wire [15:0] iffcq13pinrsrvdas;
wire [6:0]  iffcq13txsequence;
wire [1:0]  iffcq13rxdatavalid;
wire [1:0]  iffcq13rxpowerdown;
wire [1:0]  iffcq13rxresetmode;
wire [1:0]  iffcq13txbufstatus;
wire [1:0]  iffcq13txpowerdown;
wire [1:0]  iffcq13txresetmode;
wire [2:0]  iffcq13rxbufstatus;
wire [3:0]  iffcq13bufgtcemask;
wire [4:0]  iffcq13stepsizeppm;
wire [1:0]  iffcq13rxstartofseq;
wire [3:0]  iffcq13bufgtrstmask;
wire [1:0]  iffcq13rxheadervalid;
wire [2:0]  iffcq13txpmaresetmask;
wire [4:0]  iffcq13rxpcsresetmask;
wire [6:0]  iffcq13rxpmaresetmask;
wire [1:0]  iffcq13rxdapiresetmask;
wire [1:0]  iffcq13txdapiresetmask;
wire [1:0]  iffcq13rxchicoresetmask;
wire [1:0]  iffcq13txchicoresetmask;
wire [7:0]  iffcq13rxethernetstatout;

wire iffcq20enppm;
wire iffcq20perstb;
wire iffcq20bufgtce;
wire iffcq20cdrhold;
wire iffcq20cdrlock;
wire iffcq20dmonclk;
wire iffcq20rxlpmen;
wire iffcq20rxpkdet;
wire iffcq20rxqpien;
wire iffcq20rxslide;
wire iffcq20rxvalid;
wire iffcq20tstclk0;
wire iffcq20tstclk1;
wire iffcq20txswing;
wire iffcq20bufgtrst;
wire iffcq20cdrovren;
wire iffcq20cfokdone;
wire iffcq20iloreset;
wire iffcq20phyready;
wire iffcq20rxlatclk;
wire iffcq20rxusrclk;
wire iffcq20rxusrrdy;
wire iffcq20txcomsas;
wire iffcq20txlatclk;
wire iffcq20txusrclk;
wire iffcq20txusrrdy;
wire iffcq20bsrserial;
wire iffcq20cdrfreqos;
wire iffcq20cdrstepsq;
wire iffcq20cdrstepsx;
wire iffcq20comsasdet;
wire iffcq20gtrxreset;
wire iffcq20gttxreset;
wire iffcq20phystatus;
wire iffcq20rxprbserr;
wire iffcq20rxqpisenn;
wire iffcq20rxqpisenp;
wire iffcq20txcominit;
wire iffcq20txcomwake;
wire iffcq20txdccdone;
wire iffcq20txinhibit;
wire iffcq20txqpisenn;
wire iffcq20txqpisenp;
wire iffcq20aptexthold;
wire iffcq20cdrbmcdreq;
wire iffcq20cdrphreset;
wire iffcq20cdrstepdir;
wire iffcq20cominitdet;
wire iffcq20comwakedet;
wire iffcq20rxcommadet;
wire iffcq20rxelecidle;
wire iffcq20rxoobreset;
wire iffcq20rxpolarity;
wire iffcq20rxsliderdy;
wire iffcq20rxslipdone;
wire iffcq20rxsyncdone;
wire iffcq20txelecidle;
wire iffcq20txpolarity;
wire iffcq20txserpwrdn;
wire iffcq20txsyncdone;
wire iffcq20aptoverwren;
wire iffcq20cdrincpctrl;
wire iffcq20ckpinrsrvd0;
wire iffcq20ckpinrsrvd1;
wire iffcq20cssdstopclk;
wire iffcq20rxcdrphdone;
wire iffcq20rxdapireset;
wire iffcq20rxoutpcsclk;
wire iffcq20rxresetdone;
wire iffcq20rxsyncallin;
wire iffcq20txcomfinish;
wire iffcq20txdapireset;
wire iffcq20txoneszeros;
wire iffcq20txoutpcsclk;
wire iffcq20txqpibiasen;
wire iffcq20txqpiweakpu;
wire iffcq20txresetdone;
wire iffcq20txsyncallin;
wire iffcq20eyescanreset;
wire iffcq20hsdppcsreset;
wire iffcq20iloresetdone;
wire iffcq20iloresetmask;
wire iffcq20rxeqtraining;
wire iffcq20rxphdlyreset;
wire iffcq20rxprbslocked;
wire iffcq20txphdlyreset;
wire iffcq20dmonfiforeset;
wire iffcq20rxbyterealign;
wire iffcq20rxchanbondseq;
wire iffcq20rxchanrealign;
wire iffcq20rxchisaligned;
wire iffcq20rxgearboxslip;
wire iffcq20rxmldchainreq;
wire iffcq20rxtermination;
wire iffcq20txmldchainreq;
wire iffcq20txswingoutlow;
wire iffcq20eyescantrigger;
wire iffcq20resetexception;
wire iffcq20rxmldchaindone;
wire iffcq20rxphasealignpd;
wire iffcq20rxpmaresetdone;
wire iffcq20rxprbscntreset;
wire iffcq20rxprogdivreset;
wire iffcq20tcoclkfsmfrout;
wire iffcq20txchicooutrsvd;
wire iffcq20txmldchaindone;
wire iffcq20txpcsresetmask;
wire iffcq20txphasealignpd;
wire iffcq20txpmaresetdone;
wire iffcq20txprbsforceerr;
wire iffcq20txprogdivreset;
wire iffcq20txswingouthigh;
wire iffcq20rxbyteisaligned;
wire iffcq20rxdapicodereset;
wire iffcq20rxdapiresetdone;
wire iffcq20rxdelayalignerr;
wire iffcq20rxdelayalignreq;
wire iffcq20rxfinealigndone;
wire iffcq20rxphasealignerr;
wire iffcq20rxphasealignreq;
wire iffcq20txdapicodereset;
wire iffcq20txdapiresetdone;
wire iffcq20txdelayalignerr;
wire iffcq20txdelayalignreq;
wire iffcq20txphasealignerr;
wire iffcq20txphasealignreq;
wire iffcq20txtxpicodereset;
wire iffcq20eyescandataerror;
wire iffcq20rxdapicodeovrden;
wire iffcq20rxmlfinealignreq;
wire iffcq20rxphasealigndone;
wire iffcq20txdapicodeovrden;
wire iffcq20txphasealigndone;
wire iffcq20txtxpicodeovrden;
wire iffcq20xpipe5pipelineen;
wire iffcq20rxphasesetinitreq;
wire iffcq20txpausedelayalign;
wire iffcq20txphasesetinitreq;
wire iffcq20rxphasesetinitdone;
wire iffcq20rxphaseshift180req;
wire iffcq20rxprogdivresetdone;
wire iffcq20rxsimplexphystatus;
wire iffcq20txdetectrxloopback;
wire iffcq20txphasesetinitdone;
wire iffcq20txphaseshift180req;
wire iffcq20txprogdivresetdone;
wire iffcq20txsimplexphystatus;
wire iffcq20rxphaseshift180done;
wire iffcq20txphaseshift180done;
wire iffcq20phyesmadaptationsave;
wire iffcq20rxdelayalignprogress;
wire iffcq20txdelayalignprogress;
wire iffcq20rxphasedelayresetdone;
wire iffcq20txphasedelayresetdone;
wire iffcq20txethernetstattxlocalfault;

wire [7:0]  iffcq20rxrate;
wire [7:0]  iffcq20txrate;
wire[127:0] iffcq20rxdata;
wire[127:0] iffcq20txdata;
wire [15:0] iffcq20rxctrl0;
wire [15:0] iffcq20rxctrl1;
wire [15:0] iffcq20txctrl0;
wire [15:0] iffcq20txctrl1;
wire [31:0] iffcq20dmonout;
wire [7:0]  iffcq20rxctrl2;
wire [7:0]  iffcq20rxctrl3;
wire [7:0]  iffcq20txctrl2;
wire [1:0]  iffcq20txdeemph;
wire [11:0] iffcq20bufgtdiv;
wire [15:0] iffcq20pinrsrvd;
wire [2:0]  iffcq20loopback;
wire [2:0]  iffcq20rxstatus;
wire [2:0]  iffcq20txmargin;
wire [4:0]  iffcq20txdrvamp;
wire [4:0]  iffcq20txemppos;
wire [4:0]  iffcq20txemppre;
wire [5:0]  iffcq20rxheader;
wire [5:0]  iffcq20txheader;
wire [1:0]  iffcq20refclkpma;
wire [15:0] iffcq20pcsrsvdin;
wire [3:0]  iffcq20rxprbssel;
wire [3:0]  iffcq20txprbssel;
wire [4:0]  iffcq20rxchbondi;
wire [4:0]  iffcq20rxchbondo;
wire [6:0]  iffcq20txempmain;
wire [1:0]  iffcq20rxckcorcnt;
wire [15:0] iffcq20pcsrsvdout;
wire [15:0] iffcq20pinrsrvdas;
wire [6:0]  iffcq20txsequence;
wire [1:0]  iffcq20rxdatavalid;
wire [1:0]  iffcq20rxpowerdown;
wire [1:0]  iffcq20rxresetmode;
wire [1:0]  iffcq20txbufstatus;
wire [1:0]  iffcq20txpowerdown;
wire [1:0]  iffcq20txresetmode;
wire [2:0]  iffcq20rxbufstatus;
wire [3:0]  iffcq20bufgtcemask;
wire [4:0]  iffcq20stepsizeppm;
wire [1:0]  iffcq20rxstartofseq;
wire [3:0]  iffcq20bufgtrstmask;
wire [1:0]  iffcq20rxheadervalid;
wire [2:0]  iffcq20txpmaresetmask;
wire [4:0]  iffcq20rxpcsresetmask;
wire [6:0]  iffcq20rxpmaresetmask;
wire [1:0]  iffcq20rxdapiresetmask;
wire [1:0]  iffcq20txdapiresetmask;
wire [1:0]  iffcq20rxchicoresetmask;
wire [1:0]  iffcq20txchicoresetmask;
wire [7:0]  iffcq20rxethernetstatout;

wire iffcq21enppm;
wire iffcq21perstb;
wire iffcq21bufgtce;
wire iffcq21cdrhold;
wire iffcq21cdrlock;
wire iffcq21dmonclk;
wire iffcq21rxlpmen;
wire iffcq21rxpkdet;
wire iffcq21rxqpien;
wire iffcq21rxslide;
wire iffcq21rxvalid;
wire iffcq21tstclk0;
wire iffcq21tstclk1;
wire iffcq21txswing;
wire iffcq21bufgtrst;
wire iffcq21cdrovren;
wire iffcq21cfokdone;
wire iffcq21iloreset;
wire iffcq21phyready;
wire iffcq21rxlatclk;
wire iffcq21rxusrclk;
wire iffcq21rxusrrdy;
wire iffcq21txcomsas;
wire iffcq21txlatclk;
wire iffcq21txusrclk;
wire iffcq21txusrrdy;
wire iffcq21bsrserial;
wire iffcq21cdrfreqos;
wire iffcq21cdrstepsq;
wire iffcq21cdrstepsx;
wire iffcq21comsasdet;
wire iffcq21gtrxreset;
wire iffcq21gttxreset;
wire iffcq21phystatus;
wire iffcq21rxprbserr;
wire iffcq21rxqpisenn;
wire iffcq21rxqpisenp;
wire iffcq21txcominit;
wire iffcq21txcomwake;
wire iffcq21txdccdone;
wire iffcq21txinhibit;
wire iffcq21txqpisenn;
wire iffcq21txqpisenp;
wire iffcq21aptexthold;
wire iffcq21cdrbmcdreq;
wire iffcq21cdrphreset;
wire iffcq21cdrstepdir;
wire iffcq21cominitdet;
wire iffcq21comwakedet;
wire iffcq21rxcommadet;
wire iffcq21rxelecidle;
wire iffcq21rxoobreset;
wire iffcq21rxpolarity;
wire iffcq21rxsliderdy;
wire iffcq21rxslipdone;
wire iffcq21rxsyncdone;
wire iffcq21txelecidle;
wire iffcq21txpolarity;
wire iffcq21txserpwrdn;
wire iffcq21txsyncdone;
wire iffcq21aptoverwren;
wire iffcq21cdrincpctrl;
wire iffcq21ckpinrsrvd0;
wire iffcq21ckpinrsrvd1;
wire iffcq21cssdstopclk;
wire iffcq21rxcdrphdone;
wire iffcq21rxdapireset;
wire iffcq21rxoutpcsclk;
wire iffcq21rxresetdone;
wire iffcq21rxsyncallin;
wire iffcq21txcomfinish;
wire iffcq21txdapireset;
wire iffcq21txoneszeros;
wire iffcq21txoutpcsclk;
wire iffcq21txqpibiasen;
wire iffcq21txqpiweakpu;
wire iffcq21txresetdone;
wire iffcq21txsyncallin;
wire iffcq21eyescanreset;
wire iffcq21hsdppcsreset;
wire iffcq21iloresetdone;
wire iffcq21iloresetmask;
wire iffcq21rxeqtraining;
wire iffcq21rxphdlyreset;
wire iffcq21rxprbslocked;
wire iffcq21txphdlyreset;
wire iffcq21dmonfiforeset;
wire iffcq21rxbyterealign;
wire iffcq21rxchanbondseq;
wire iffcq21rxchanrealign;
wire iffcq21rxchisaligned;
wire iffcq21rxgearboxslip;
wire iffcq21rxmldchainreq;
wire iffcq21rxtermination;
wire iffcq21txmldchainreq;
wire iffcq21txswingoutlow;
wire iffcq21eyescantrigger;
wire iffcq21resetexception;
wire iffcq21rxmldchaindone;
wire iffcq21rxphasealignpd;
wire iffcq21rxpmaresetdone;
wire iffcq21rxprbscntreset;
wire iffcq21rxprogdivreset;
wire iffcq21tcoclkfsmfrout;
wire iffcq21txchicooutrsvd;
wire iffcq21txmldchaindone;
wire iffcq21txpcsresetmask;
wire iffcq21txphasealignpd;
wire iffcq21txpmaresetdone;
wire iffcq21txprbsforceerr;
wire iffcq21txprogdivreset;
wire iffcq21txswingouthigh;
wire iffcq21rxbyteisaligned;
wire iffcq21rxdapicodereset;
wire iffcq21rxdapiresetdone;
wire iffcq21rxdelayalignerr;
wire iffcq21rxdelayalignreq;
wire iffcq21rxfinealigndone;
wire iffcq21rxphasealignerr;
wire iffcq21rxphasealignreq;
wire iffcq21txdapicodereset;
wire iffcq21txdapiresetdone;
wire iffcq21txdelayalignerr;
wire iffcq21txdelayalignreq;
wire iffcq21txphasealignerr;
wire iffcq21txphasealignreq;
wire iffcq21txtxpicodereset;
wire iffcq21eyescandataerror;
wire iffcq21rxdapicodeovrden;
wire iffcq21rxmlfinealignreq;
wire iffcq21rxphasealigndone;
wire iffcq21txdapicodeovrden;
wire iffcq21txphasealigndone;
wire iffcq21txtxpicodeovrden;
wire iffcq21xpipe5pipelineen;
wire iffcq21rxphasesetinitreq;
wire iffcq21txpausedelayalign;
wire iffcq21txphasesetinitreq;
wire iffcq21rxphasesetinitdone;
wire iffcq21rxphaseshift180req;
wire iffcq21rxprogdivresetdone;
wire iffcq21rxsimplexphystatus;
wire iffcq21txdetectrxloopback;
wire iffcq21txphasesetinitdone;
wire iffcq21txphaseshift180req;
wire iffcq21txprogdivresetdone;
wire iffcq21txsimplexphystatus;
wire iffcq21rxphaseshift180done;
wire iffcq21txphaseshift180done;
wire iffcq21phyesmadaptationsave;
wire iffcq21rxdelayalignprogress;
wire iffcq21txdelayalignprogress;
wire iffcq21rxphasedelayresetdone;
wire iffcq21txphasedelayresetdone;
wire iffcq21txethernetstattxlocalfault;

wire [7:0]  iffcq21rxrate;
wire [7:0]  iffcq21txrate;
wire[127:0] iffcq21rxdata;
wire[127:0] iffcq21txdata;
wire [15:0] iffcq21rxctrl0;
wire [15:0] iffcq21rxctrl1;
wire [15:0] iffcq21txctrl0;
wire [15:0] iffcq21txctrl1;
wire [31:0] iffcq21dmonout;
wire [7:0]  iffcq21rxctrl2;
wire [7:0]  iffcq21rxctrl3;
wire [7:0]  iffcq21txctrl2;
wire [1:0]  iffcq21txdeemph;
wire [11:0] iffcq21bufgtdiv;
wire [15:0] iffcq21pinrsrvd;
wire [2:0]  iffcq21loopback;
wire [2:0]  iffcq21rxstatus;
wire [2:0]  iffcq21txmargin;
wire [4:0]  iffcq21txdrvamp;
wire [4:0]  iffcq21txemppos;
wire [4:0]  iffcq21txemppre;
wire [5:0]  iffcq21rxheader;
wire [5:0]  iffcq21txheader;
wire [1:0]  iffcq21refclkpma;
wire [15:0] iffcq21pcsrsvdin;
wire [3:0]  iffcq21rxprbssel;
wire [3:0]  iffcq21txprbssel;
wire [4:0]  iffcq21rxchbondi;
wire [4:0]  iffcq21rxchbondo;
wire [6:0]  iffcq21txempmain;
wire [1:0]  iffcq21rxckcorcnt;
wire [15:0] iffcq21pcsrsvdout;
wire [15:0] iffcq21pinrsrvdas;
wire [6:0]  iffcq21txsequence;
wire [1:0]  iffcq21rxdatavalid;
wire [1:0]  iffcq21rxpowerdown;
wire [1:0]  iffcq21rxresetmode;
wire [1:0]  iffcq21txbufstatus;
wire [1:0]  iffcq21txpowerdown;
wire [1:0]  iffcq21txresetmode;
wire [2:0]  iffcq21rxbufstatus;
wire [3:0]  iffcq21bufgtcemask;
wire [4:0]  iffcq21stepsizeppm;
wire [1:0]  iffcq21rxstartofseq;
wire [3:0]  iffcq21bufgtrstmask;
wire [1:0]  iffcq21rxheadervalid;
wire [2:0]  iffcq21txpmaresetmask;
wire [4:0]  iffcq21rxpcsresetmask;
wire [6:0]  iffcq21rxpmaresetmask;
wire [1:0]  iffcq21rxdapiresetmask;
wire [1:0]  iffcq21txdapiresetmask;
wire [1:0]  iffcq21rxchicoresetmask;
wire [1:0]  iffcq21txchicoresetmask;
wire [7:0]  iffcq21rxethernetstatout;

wire iffcq22enppm;
wire iffcq22perstb;
wire iffcq22bufgtce;
wire iffcq22cdrhold;
wire iffcq22cdrlock;
wire iffcq22dmonclk;
wire iffcq22rxlpmen;
wire iffcq22rxpkdet;
wire iffcq22rxqpien;
wire iffcq22rxslide;
wire iffcq22rxvalid;
wire iffcq22tstclk0;
wire iffcq22tstclk1;
wire iffcq22txswing;
wire iffcq22bufgtrst;
wire iffcq22cdrovren;
wire iffcq22cfokdone;
wire iffcq22iloreset;
wire iffcq22phyready;
wire iffcq22rxlatclk;
wire iffcq22rxusrclk;
wire iffcq22rxusrrdy;
wire iffcq22txcomsas;
wire iffcq22txlatclk;
wire iffcq22txusrclk;
wire iffcq22txusrrdy;
wire iffcq22bsrserial;
wire iffcq22cdrfreqos;
wire iffcq22cdrstepsq;
wire iffcq22cdrstepsx;
wire iffcq22comsasdet;
wire iffcq22gtrxreset;
wire iffcq22gttxreset;
wire iffcq22phystatus;
wire iffcq22rxprbserr;
wire iffcq22rxqpisenn;
wire iffcq22rxqpisenp;
wire iffcq22txcominit;
wire iffcq22txcomwake;
wire iffcq22txdccdone;
wire iffcq22txinhibit;
wire iffcq22txqpisenn;
wire iffcq22txqpisenp;
wire iffcq22aptexthold;
wire iffcq22cdrbmcdreq;
wire iffcq22cdrphreset;
wire iffcq22cdrstepdir;
wire iffcq22cominitdet;
wire iffcq22comwakedet;
wire iffcq22rxcommadet;
wire iffcq22rxelecidle;
wire iffcq22rxoobreset;
wire iffcq22rxpolarity;
wire iffcq22rxsliderdy;
wire iffcq22rxslipdone;
wire iffcq22rxsyncdone;
wire iffcq22txelecidle;
wire iffcq22txpolarity;
wire iffcq22txserpwrdn;
wire iffcq22txsyncdone;
wire iffcq22aptoverwren;
wire iffcq22cdrincpctrl;
wire iffcq22ckpinrsrvd0;
wire iffcq22ckpinrsrvd1;
wire iffcq22cssdstopclk;
wire iffcq22rxcdrphdone;
wire iffcq22rxdapireset;
wire iffcq22rxoutpcsclk;
wire iffcq22rxresetdone;
wire iffcq22rxsyncallin;
wire iffcq22txcomfinish;
wire iffcq22txdapireset;
wire iffcq22txoneszeros;
wire iffcq22txoutpcsclk;
wire iffcq22txqpibiasen;
wire iffcq22txqpiweakpu;
wire iffcq22txresetdone;
wire iffcq22txsyncallin;
wire iffcq22eyescanreset;
wire iffcq22hsdppcsreset;
wire iffcq22iloresetdone;
wire iffcq22iloresetmask;
wire iffcq22rxeqtraining;
wire iffcq22rxphdlyreset;
wire iffcq22rxprbslocked;
wire iffcq22txphdlyreset;
wire iffcq22dmonfiforeset;
wire iffcq22rxbyterealign;
wire iffcq22rxchanbondseq;
wire iffcq22rxchanrealign;
wire iffcq22rxchisaligned;
wire iffcq22rxgearboxslip;
wire iffcq22rxmldchainreq;
wire iffcq22rxtermination;
wire iffcq22txmldchainreq;
wire iffcq22txswingoutlow;
wire iffcq22eyescantrigger;
wire iffcq22resetexception;
wire iffcq22rxmldchaindone;
wire iffcq22rxphasealignpd;
wire iffcq22rxpmaresetdone;
wire iffcq22rxprbscntreset;
wire iffcq22rxprogdivreset;
wire iffcq22tcoclkfsmfrout;
wire iffcq22txchicooutrsvd;
wire iffcq22txmldchaindone;
wire iffcq22txpcsresetmask;
wire iffcq22txphasealignpd;
wire iffcq22txpmaresetdone;
wire iffcq22txprbsforceerr;
wire iffcq22txprogdivreset;
wire iffcq22txswingouthigh;
wire iffcq22rxbyteisaligned;
wire iffcq22rxdapicodereset;
wire iffcq22rxdapiresetdone;
wire iffcq22rxdelayalignerr;
wire iffcq22rxdelayalignreq;
wire iffcq22rxfinealigndone;
wire iffcq22rxphasealignerr;
wire iffcq22rxphasealignreq;
wire iffcq22txdapicodereset;
wire iffcq22txdapiresetdone;
wire iffcq22txdelayalignerr;
wire iffcq22txdelayalignreq;
wire iffcq22txphasealignerr;
wire iffcq22txphasealignreq;
wire iffcq22txtxpicodereset;
wire iffcq22eyescandataerror;
wire iffcq22rxdapicodeovrden;
wire iffcq22rxmlfinealignreq;
wire iffcq22rxphasealigndone;
wire iffcq22txdapicodeovrden;
wire iffcq22txphasealigndone;
wire iffcq22txtxpicodeovrden;
wire iffcq22xpipe5pipelineen;
wire iffcq22rxphasesetinitreq;
wire iffcq22txpausedelayalign;
wire iffcq22txphasesetinitreq;
wire iffcq22rxphasesetinitdone;
wire iffcq22rxphaseshift180req;
wire iffcq22rxprogdivresetdone;
wire iffcq22rxsimplexphystatus;
wire iffcq22txdetectrxloopback;
wire iffcq22txphasesetinitdone;
wire iffcq22txphaseshift180req;
wire iffcq22txprogdivresetdone;
wire iffcq22txsimplexphystatus;
wire iffcq22rxphaseshift180done;
wire iffcq22txphaseshift180done;
wire iffcq22phyesmadaptationsave;
wire iffcq22rxdelayalignprogress;
wire iffcq22txdelayalignprogress;
wire iffcq22rxphasedelayresetdone;
wire iffcq22txphasedelayresetdone;
wire iffcq22txethernetstattxlocalfault;

wire [7:0]  iffcq22rxrate;
wire [7:0]  iffcq22txrate;
wire[127:0] iffcq22rxdata;
wire[127:0] iffcq22txdata;
wire [15:0] iffcq22rxctrl0;
wire [15:0] iffcq22rxctrl1;
wire [15:0] iffcq22txctrl0;
wire [15:0] iffcq22txctrl1;
wire [31:0] iffcq22dmonout;
wire [7:0]  iffcq22rxctrl2;
wire [7:0]  iffcq22rxctrl3;
wire [7:0]  iffcq22txctrl2;
wire [1:0]  iffcq22txdeemph;
wire [11:0] iffcq22bufgtdiv;
wire [15:0] iffcq22pinrsrvd;
wire [2:0]  iffcq22loopback;
wire [2:0]  iffcq22rxstatus;
wire [2:0]  iffcq22txmargin;
wire [4:0]  iffcq22txdrvamp;
wire [4:0]  iffcq22txemppos;
wire [4:0]  iffcq22txemppre;
wire [5:0]  iffcq22rxheader;
wire [5:0]  iffcq22txheader;
wire [1:0]  iffcq22refclkpma;
wire [15:0] iffcq22pcsrsvdin;
wire [3:0]  iffcq22rxprbssel;
wire [3:0]  iffcq22txprbssel;
wire [4:0]  iffcq22rxchbondi;
wire [4:0]  iffcq22rxchbondo;
wire [6:0]  iffcq22txempmain;
wire [1:0]  iffcq22rxckcorcnt;
wire [15:0] iffcq22pcsrsvdout;
wire [15:0] iffcq22pinrsrvdas;
wire [6:0]  iffcq22txsequence;
wire [1:0]  iffcq22rxdatavalid;
wire [1:0]  iffcq22rxpowerdown;
wire [1:0]  iffcq22rxresetmode;
wire [1:0]  iffcq22txbufstatus;
wire [1:0]  iffcq22txpowerdown;
wire [1:0]  iffcq22txresetmode;
wire [2:0]  iffcq22rxbufstatus;
wire [3:0]  iffcq22bufgtcemask;
wire [4:0]  iffcq22stepsizeppm;
wire [1:0]  iffcq22rxstartofseq;
wire [3:0]  iffcq22bufgtrstmask;
wire [1:0]  iffcq22rxheadervalid;
wire [2:0]  iffcq22txpmaresetmask;
wire [4:0]  iffcq22rxpcsresetmask;
wire [6:0]  iffcq22rxpmaresetmask;
wire [1:0]  iffcq22rxdapiresetmask;
wire [1:0]  iffcq22txdapiresetmask;
wire [1:0]  iffcq22rxchicoresetmask;
wire [1:0]  iffcq22txchicoresetmask;
wire [7:0]  iffcq22rxethernetstatout;

wire iffcq23enppm;
wire iffcq23perstb;
wire iffcq23bufgtce;
wire iffcq23cdrhold;
wire iffcq23cdrlock;
wire iffcq23dmonclk;
wire iffcq23rxlpmen;
wire iffcq23rxpkdet;
wire iffcq23rxqpien;
wire iffcq23rxslide;
wire iffcq23rxvalid;
wire iffcq23tstclk0;
wire iffcq23tstclk1;
wire iffcq23txswing;
wire iffcq23bufgtrst;
wire iffcq23cdrovren;
wire iffcq23cfokdone;
wire iffcq23iloreset;
wire iffcq23phyready;
wire iffcq23rxlatclk;
wire iffcq23rxusrclk;
wire iffcq23rxusrrdy;
wire iffcq23txcomsas;
wire iffcq23txlatclk;
wire iffcq23txusrclk;
wire iffcq23txusrrdy;
wire iffcq23bsrserial;
wire iffcq23cdrfreqos;
wire iffcq23cdrstepsq;
wire iffcq23cdrstepsx;
wire iffcq23comsasdet;
wire iffcq23gtrxreset;
wire iffcq23gttxreset;
wire iffcq23phystatus;
wire iffcq23rxprbserr;
wire iffcq23rxqpisenn;
wire iffcq23rxqpisenp;
wire iffcq23txcominit;
wire iffcq23txcomwake;
wire iffcq23txdccdone;
wire iffcq23txinhibit;
wire iffcq23txqpisenn;
wire iffcq23txqpisenp;
wire iffcq23aptexthold;
wire iffcq23cdrbmcdreq;
wire iffcq23cdrphreset;
wire iffcq23cdrstepdir;
wire iffcq23cominitdet;
wire iffcq23comwakedet;
wire iffcq23rxcommadet;
wire iffcq23rxelecidle;
wire iffcq23rxoobreset;
wire iffcq23rxpolarity;
wire iffcq23rxsliderdy;
wire iffcq23rxslipdone;
wire iffcq23rxsyncdone;
wire iffcq23txelecidle;
wire iffcq23txpolarity;
wire iffcq23txserpwrdn;
wire iffcq23txsyncdone;
wire iffcq23aptoverwren;
wire iffcq23cdrincpctrl;
wire iffcq23ckpinrsrvd0;
wire iffcq23ckpinrsrvd1;
wire iffcq23cssdstopclk;
wire iffcq23rxcdrphdone;
wire iffcq23rxdapireset;
wire iffcq23rxoutpcsclk;
wire iffcq23rxresetdone;
wire iffcq23rxsyncallin;
wire iffcq23txcomfinish;
wire iffcq23txdapireset;
wire iffcq23txoneszeros;
wire iffcq23txoutpcsclk;
wire iffcq23txqpibiasen;
wire iffcq23txqpiweakpu;
wire iffcq23txresetdone;
wire iffcq23txsyncallin;
wire iffcq23eyescanreset;
wire iffcq23hsdppcsreset;
wire iffcq23iloresetdone;
wire iffcq23iloresetmask;
wire iffcq23rxeqtraining;
wire iffcq23rxphdlyreset;
wire iffcq23rxprbslocked;
wire iffcq23txphdlyreset;
wire iffcq23dmonfiforeset;
wire iffcq23rxbyterealign;
wire iffcq23rxchanbondseq;
wire iffcq23rxchanrealign;
wire iffcq23rxchisaligned;
wire iffcq23rxgearboxslip;
wire iffcq23rxmldchainreq;
wire iffcq23rxtermination;
wire iffcq23txmldchainreq;
wire iffcq23txswingoutlow;
wire iffcq23eyescantrigger;
wire iffcq23resetexception;
wire iffcq23rxmldchaindone;
wire iffcq23rxphasealignpd;
wire iffcq23rxpmaresetdone;
wire iffcq23rxprbscntreset;
wire iffcq23rxprogdivreset;
wire iffcq23tcoclkfsmfrout;
wire iffcq23txchicooutrsvd;
wire iffcq23txmldchaindone;
wire iffcq23txpcsresetmask;
wire iffcq23txphasealignpd;
wire iffcq23txpmaresetdone;
wire iffcq23txprbsforceerr;
wire iffcq23txprogdivreset;
wire iffcq23txswingouthigh;
wire iffcq23rxbyteisaligned;
wire iffcq23rxdapicodereset;
wire iffcq23rxdapiresetdone;
wire iffcq23rxdelayalignerr;
wire iffcq23rxdelayalignreq;
wire iffcq23rxfinealigndone;
wire iffcq23rxphasealignerr;
wire iffcq23rxphasealignreq;
wire iffcq23txdapicodereset;
wire iffcq23txdapiresetdone;
wire iffcq23txdelayalignerr;
wire iffcq23txdelayalignreq;
wire iffcq23txphasealignerr;
wire iffcq23txphasealignreq;
wire iffcq23txtxpicodereset;
wire iffcq23eyescandataerror;
wire iffcq23rxdapicodeovrden;
wire iffcq23rxmlfinealignreq;
wire iffcq23rxphasealigndone;
wire iffcq23txdapicodeovrden;
wire iffcq23txphasealigndone;
wire iffcq23txtxpicodeovrden;
wire iffcq23xpipe5pipelineen;
wire iffcq23rxphasesetinitreq;
wire iffcq23txpausedelayalign;
wire iffcq23txphasesetinitreq;
wire iffcq23rxphasesetinitdone;
wire iffcq23rxphaseshift180req;
wire iffcq23rxprogdivresetdone;
wire iffcq23rxsimplexphystatus;
wire iffcq23txdetectrxloopback;
wire iffcq23txphasesetinitdone;
wire iffcq23txphaseshift180req;
wire iffcq23txprogdivresetdone;
wire iffcq23txsimplexphystatus;
wire iffcq23rxphaseshift180done;
wire iffcq23txphaseshift180done;
wire iffcq23phyesmadaptationsave;
wire iffcq23rxdelayalignprogress;
wire iffcq23txdelayalignprogress;
wire iffcq23rxphasedelayresetdone;
wire iffcq23txphasedelayresetdone;
wire iffcq23txethernetstattxlocalfault;

wire [7:0]  iffcq23rxrate;
wire [7:0]  iffcq23txrate;
wire[127:0] iffcq23rxdata;
wire[127:0] iffcq23txdata;
wire [15:0] iffcq23rxctrl0;
wire [15:0] iffcq23rxctrl1;
wire [15:0] iffcq23txctrl0;
wire [15:0] iffcq23txctrl1;
wire [31:0] iffcq23dmonout;
wire [7:0]  iffcq23rxctrl2;
wire [7:0]  iffcq23rxctrl3;
wire [7:0]  iffcq23txctrl2;
wire [1:0]  iffcq23txdeemph;
wire [11:0] iffcq23bufgtdiv;
wire [15:0] iffcq23pinrsrvd;
wire [2:0]  iffcq23loopback;
wire [2:0]  iffcq23rxstatus;
wire [2:0]  iffcq23txmargin;
wire [4:0]  iffcq23txdrvamp;
wire [4:0]  iffcq23txemppos;
wire [4:0]  iffcq23txemppre;
wire [5:0]  iffcq23rxheader;
wire [5:0]  iffcq23txheader;
wire [1:0]  iffcq23refclkpma;
wire [15:0] iffcq23pcsrsvdin;
wire [3:0]  iffcq23rxprbssel;
wire [3:0]  iffcq23txprbssel;
wire [4:0]  iffcq23rxchbondi;
wire [4:0]  iffcq23rxchbondo;
wire [6:0]  iffcq23txempmain;
wire [1:0]  iffcq23rxckcorcnt;
wire [15:0] iffcq23pcsrsvdout;
wire [15:0] iffcq23pinrsrvdas;
wire [6:0]  iffcq23txsequence;
wire [1:0]  iffcq23rxdatavalid;
wire [1:0]  iffcq23rxpowerdown;
wire [1:0]  iffcq23rxresetmode;
wire [1:0]  iffcq23txbufstatus;
wire [1:0]  iffcq23txpowerdown;
wire [1:0]  iffcq23txresetmode;
wire [2:0]  iffcq23rxbufstatus;
wire [3:0]  iffcq23bufgtcemask;
wire [4:0]  iffcq23stepsizeppm;
wire [1:0]  iffcq23rxstartofseq;
wire [3:0]  iffcq23bufgtrstmask;
wire [1:0]  iffcq23rxheadervalid;
wire [2:0]  iffcq23txpmaresetmask;
wire [4:0]  iffcq23rxpcsresetmask;
wire [6:0]  iffcq23rxpmaresetmask;
wire [1:0]  iffcq23rxdapiresetmask;
wire [1:0]  iffcq23txdapiresetmask;
wire [1:0]  iffcq23rxchicoresetmask;
wire [1:0]  iffcq23txchicoresetmask;
wire [7:0]  iffcq23rxethernetstatout;

wire iffcq30enppm;
wire iffcq30perstb;
wire iffcq30bufgtce;
wire iffcq30cdrhold;
wire iffcq30cdrlock;
wire iffcq30dmonclk;
wire iffcq30rxlpmen;
wire iffcq30rxpkdet;
wire iffcq30rxqpien;
wire iffcq30rxslide;
wire iffcq30rxvalid;
wire iffcq30tstclk0;
wire iffcq30tstclk1;
wire iffcq30txswing;
wire iffcq30bufgtrst;
wire iffcq30cdrovren;
wire iffcq30cfokdone;
wire iffcq30iloreset;
wire iffcq30phyready;
wire iffcq30rxlatclk;
wire iffcq30rxusrclk;
wire iffcq30rxusrrdy;
wire iffcq30txcomsas;
wire iffcq30txlatclk;
wire iffcq30txusrclk;
wire iffcq30txusrrdy;
wire iffcq30bsrserial;
wire iffcq30cdrfreqos;
wire iffcq30cdrstepsq;
wire iffcq30cdrstepsx;
wire iffcq30comsasdet;
wire iffcq30gtrxreset;
wire iffcq30gttxreset;
wire iffcq30phystatus;
wire iffcq30rxprbserr;
wire iffcq30rxqpisenn;
wire iffcq30rxqpisenp;
wire iffcq30txcominit;
wire iffcq30txcomwake;
wire iffcq30txdccdone;
wire iffcq30txinhibit;
wire iffcq30txqpisenn;
wire iffcq30txqpisenp;
wire iffcq30aptexthold;
wire iffcq30cdrbmcdreq;
wire iffcq30cdrphreset;
wire iffcq30cdrstepdir;
wire iffcq30cominitdet;
wire iffcq30comwakedet;
wire iffcq30rxcommadet;
wire iffcq30rxelecidle;
wire iffcq30rxoobreset;
wire iffcq30rxpolarity;
wire iffcq30rxsliderdy;
wire iffcq30rxslipdone;
wire iffcq30rxsyncdone;
wire iffcq30txelecidle;
wire iffcq30txpolarity;
wire iffcq30txserpwrdn;
wire iffcq30txsyncdone;
wire iffcq30aptoverwren;
wire iffcq30cdrincpctrl;
wire iffcq30ckpinrsrvd0;
wire iffcq30ckpinrsrvd1;
wire iffcq30cssdstopclk;
wire iffcq30rxcdrphdone;
wire iffcq30rxdapireset;
wire iffcq30rxoutpcsclk;
wire iffcq30rxresetdone;
wire iffcq30rxsyncallin;
wire iffcq30txcomfinish;
wire iffcq30txdapireset;
wire iffcq30txoneszeros;
wire iffcq30txoutpcsclk;
wire iffcq30txqpibiasen;
wire iffcq30txqpiweakpu;
wire iffcq30txresetdone;
wire iffcq30txsyncallin;
wire iffcq30eyescanreset;
wire iffcq30hsdppcsreset;
wire iffcq30iloresetdone;
wire iffcq30iloresetmask;
wire iffcq30rxeqtraining;
wire iffcq30rxphdlyreset;
wire iffcq30rxprbslocked;
wire iffcq30txphdlyreset;
wire iffcq30dmonfiforeset;
wire iffcq30rxbyterealign;
wire iffcq30rxchanbondseq;
wire iffcq30rxchanrealign;
wire iffcq30rxchisaligned;
wire iffcq30rxgearboxslip;
wire iffcq30rxmldchainreq;
wire iffcq30rxtermination;
wire iffcq30txmldchainreq;
wire iffcq30txswingoutlow;
wire iffcq30eyescantrigger;
wire iffcq30resetexception;
wire iffcq30rxmldchaindone;
wire iffcq30rxphasealignpd;
wire iffcq30rxpmaresetdone;
wire iffcq30rxprbscntreset;
wire iffcq30rxprogdivreset;
wire iffcq30tcoclkfsmfrout;
wire iffcq30txchicooutrsvd;
wire iffcq30txmldchaindone;
wire iffcq30txpcsresetmask;
wire iffcq30txphasealignpd;
wire iffcq30txpmaresetdone;
wire iffcq30txprbsforceerr;
wire iffcq30txprogdivreset;
wire iffcq30txswingouthigh;
wire iffcq30rxbyteisaligned;
wire iffcq30rxdapicodereset;
wire iffcq30rxdapiresetdone;
wire iffcq30rxdelayalignerr;
wire iffcq30rxdelayalignreq;
wire iffcq30rxfinealigndone;
wire iffcq30rxphasealignerr;
wire iffcq30rxphasealignreq;
wire iffcq30txdapicodereset;
wire iffcq30txdapiresetdone;
wire iffcq30txdelayalignerr;
wire iffcq30txdelayalignreq;
wire iffcq30txphasealignerr;
wire iffcq30txphasealignreq;
wire iffcq30txtxpicodereset;
wire iffcq30eyescandataerror;
wire iffcq30rxdapicodeovrden;
wire iffcq30rxmlfinealignreq;
wire iffcq30rxphasealigndone;
wire iffcq30txdapicodeovrden;
wire iffcq30txphasealigndone;
wire iffcq30txtxpicodeovrden;
wire iffcq30xpipe5pipelineen;
wire iffcq30rxphasesetinitreq;
wire iffcq30txpausedelayalign;
wire iffcq30txphasesetinitreq;
wire iffcq30rxphasesetinitdone;
wire iffcq30rxphaseshift180req;
wire iffcq30rxprogdivresetdone;
wire iffcq30rxsimplexphystatus;
wire iffcq30txdetectrxloopback;
wire iffcq30txphasesetinitdone;
wire iffcq30txphaseshift180req;
wire iffcq30txprogdivresetdone;
wire iffcq30txsimplexphystatus;
wire iffcq30rxphaseshift180done;
wire iffcq30txphaseshift180done;
wire iffcq30phyesmadaptationsave;
wire iffcq30rxdelayalignprogress;
wire iffcq30txdelayalignprogress;
wire iffcq30rxphasedelayresetdone;
wire iffcq30txphasedelayresetdone;
wire iffcq30txethernetstattxlocalfault;

wire [7:0]  iffcq30rxrate;
wire [7:0]  iffcq30txrate;
wire[127:0] iffcq30rxdata;
wire[127:0] iffcq30txdata;
wire [15:0] iffcq30rxctrl0;
wire [15:0] iffcq30rxctrl1;
wire [15:0] iffcq30txctrl0;
wire [15:0] iffcq30txctrl1;
wire [31:0] iffcq30dmonout;
wire [7:0]  iffcq30rxctrl2;
wire [7:0]  iffcq30rxctrl3;
wire [7:0]  iffcq30txctrl2;
wire [1:0]  iffcq30txdeemph;
wire [11:0] iffcq30bufgtdiv;
wire [15:0] iffcq30pinrsrvd;
wire [2:0]  iffcq30loopback;
wire [2:0]  iffcq30rxstatus;
wire [2:0]  iffcq30txmargin;
wire [4:0]  iffcq30txdrvamp;
wire [4:0]  iffcq30txemppos;
wire [4:0]  iffcq30txemppre;
wire [5:0]  iffcq30rxheader;
wire [5:0]  iffcq30txheader;
wire [1:0]  iffcq30refclkpma;
wire [15:0] iffcq30pcsrsvdin;
wire [3:0]  iffcq30rxprbssel;
wire [3:0]  iffcq30txprbssel;
wire [4:0]  iffcq30rxchbondi;
wire [4:0]  iffcq30rxchbondo;
wire [6:0]  iffcq30txempmain;
wire [1:0]  iffcq30rxckcorcnt;
wire [15:0] iffcq30pcsrsvdout;
wire [15:0] iffcq30pinrsrvdas;
wire [6:0]  iffcq30txsequence;
wire [1:0]  iffcq30rxdatavalid;
wire [1:0]  iffcq30rxpowerdown;
wire [1:0]  iffcq30rxresetmode;
wire [1:0]  iffcq30txbufstatus;
wire [1:0]  iffcq30txpowerdown;
wire [1:0]  iffcq30txresetmode;
wire [2:0]  iffcq30rxbufstatus;
wire [3:0]  iffcq30bufgtcemask;
wire [4:0]  iffcq30stepsizeppm;
wire [1:0]  iffcq30rxstartofseq;
wire [3:0]  iffcq30bufgtrstmask;
wire [1:0]  iffcq30rxheadervalid;
wire [2:0]  iffcq30txpmaresetmask;
wire [4:0]  iffcq30rxpcsresetmask;
wire [6:0]  iffcq30rxpmaresetmask;
wire [1:0]  iffcq30rxdapiresetmask;
wire [1:0]  iffcq30txdapiresetmask;
wire [1:0]  iffcq30rxchicoresetmask;
wire [1:0]  iffcq30txchicoresetmask;
wire [7:0]  iffcq30rxethernetstatout;

wire iffcq31enppm;
wire iffcq31perstb;
wire iffcq31bufgtce;
wire iffcq31cdrhold;
wire iffcq31cdrlock;
wire iffcq31dmonclk;
wire iffcq31rxlpmen;
wire iffcq31rxpkdet;
wire iffcq31rxqpien;
wire iffcq31rxslide;
wire iffcq31rxvalid;
wire iffcq31tstclk0;
wire iffcq31tstclk1;
wire iffcq31txswing;
wire iffcq31bufgtrst;
wire iffcq31cdrovren;
wire iffcq31cfokdone;
wire iffcq31iloreset;
wire iffcq31phyready;
wire iffcq31rxlatclk;
wire iffcq31rxusrclk;
wire iffcq31rxusrrdy;
wire iffcq31txcomsas;
wire iffcq31txlatclk;
wire iffcq31txusrclk;
wire iffcq31txusrrdy;
wire iffcq31bsrserial;
wire iffcq31cdrfreqos;
wire iffcq31cdrstepsq;
wire iffcq31cdrstepsx;
wire iffcq31comsasdet;
wire iffcq31gtrxreset;
wire iffcq31gttxreset;
wire iffcq31phystatus;
wire iffcq31rxprbserr;
wire iffcq31rxqpisenn;
wire iffcq31rxqpisenp;
wire iffcq31txcominit;
wire iffcq31txcomwake;
wire iffcq31txdccdone;
wire iffcq31txinhibit;
wire iffcq31txqpisenn;
wire iffcq31txqpisenp;
wire iffcq31aptexthold;
wire iffcq31cdrbmcdreq;
wire iffcq31cdrphreset;
wire iffcq31cdrstepdir;
wire iffcq31cominitdet;
wire iffcq31comwakedet;
wire iffcq31rxcommadet;
wire iffcq31rxelecidle;
wire iffcq31rxoobreset;
wire iffcq31rxpolarity;
wire iffcq31rxsliderdy;
wire iffcq31rxslipdone;
wire iffcq31rxsyncdone;
wire iffcq31txelecidle;
wire iffcq31txpolarity;
wire iffcq31txserpwrdn;
wire iffcq31txsyncdone;
wire iffcq31aptoverwren;
wire iffcq31cdrincpctrl;
wire iffcq31ckpinrsrvd0;
wire iffcq31ckpinrsrvd1;
wire iffcq31cssdstopclk;
wire iffcq31rxcdrphdone;
wire iffcq31rxdapireset;
wire iffcq31rxoutpcsclk;
wire iffcq31rxresetdone;
wire iffcq31rxsyncallin;
wire iffcq31txcomfinish;
wire iffcq31txdapireset;
wire iffcq31txoneszeros;
wire iffcq31txoutpcsclk;
wire iffcq31txqpibiasen;
wire iffcq31txqpiweakpu;
wire iffcq31txresetdone;
wire iffcq31txsyncallin;
wire iffcq31eyescanreset;
wire iffcq31hsdppcsreset;
wire iffcq31iloresetdone;
wire iffcq31iloresetmask;
wire iffcq31rxeqtraining;
wire iffcq31rxphdlyreset;
wire iffcq31rxprbslocked;
wire iffcq31txphdlyreset;
wire iffcq31dmonfiforeset;
wire iffcq31rxbyterealign;
wire iffcq31rxchanbondseq;
wire iffcq31rxchanrealign;
wire iffcq31rxchisaligned;
wire iffcq31rxgearboxslip;
wire iffcq31rxmldchainreq;
wire iffcq31rxtermination;
wire iffcq31txmldchainreq;
wire iffcq31txswingoutlow;
wire iffcq31eyescantrigger;
wire iffcq31resetexception;
wire iffcq31rxmldchaindone;
wire iffcq31rxphasealignpd;
wire iffcq31rxpmaresetdone;
wire iffcq31rxprbscntreset;
wire iffcq31rxprogdivreset;
wire iffcq31tcoclkfsmfrout;
wire iffcq31txchicooutrsvd;
wire iffcq31txmldchaindone;
wire iffcq31txpcsresetmask;
wire iffcq31txphasealignpd;
wire iffcq31txpmaresetdone;
wire iffcq31txprbsforceerr;
wire iffcq31txprogdivreset;
wire iffcq31txswingouthigh;
wire iffcq31rxbyteisaligned;
wire iffcq31rxdapicodereset;
wire iffcq31rxdapiresetdone;
wire iffcq31rxdelayalignerr;
wire iffcq31rxdelayalignreq;
wire iffcq31rxfinealigndone;
wire iffcq31rxphasealignerr;
wire iffcq31rxphasealignreq;
wire iffcq31txdapicodereset;
wire iffcq31txdapiresetdone;
wire iffcq31txdelayalignerr;
wire iffcq31txdelayalignreq;
wire iffcq31txphasealignerr;
wire iffcq31txphasealignreq;
wire iffcq31txtxpicodereset;
wire iffcq31eyescandataerror;
wire iffcq31rxdapicodeovrden;
wire iffcq31rxmlfinealignreq;
wire iffcq31rxphasealigndone;
wire iffcq31txdapicodeovrden;
wire iffcq31txphasealigndone;
wire iffcq31txtxpicodeovrden;
wire iffcq31xpipe5pipelineen;
wire iffcq31rxphasesetinitreq;
wire iffcq31txpausedelayalign;
wire iffcq31txphasesetinitreq;
wire iffcq31rxphasesetinitdone;
wire iffcq31rxphaseshift180req;
wire iffcq31rxprogdivresetdone;
wire iffcq31rxsimplexphystatus;
wire iffcq31txdetectrxloopback;
wire iffcq31txphasesetinitdone;
wire iffcq31txphaseshift180req;
wire iffcq31txprogdivresetdone;
wire iffcq31txsimplexphystatus;
wire iffcq31rxphaseshift180done;
wire iffcq31txphaseshift180done;
wire iffcq31phyesmadaptationsave;
wire iffcq31rxdelayalignprogress;
wire iffcq31txdelayalignprogress;
wire iffcq31rxphasedelayresetdone;
wire iffcq31txphasedelayresetdone;
wire iffcq31txethernetstattxlocalfault;

wire [7:0]  iffcq31rxrate;
wire [7:0]  iffcq31txrate;
wire[127:0] iffcq31rxdata;
wire[127:0] iffcq31txdata;
wire [15:0] iffcq31rxctrl0;
wire [15:0] iffcq31rxctrl1;
wire [15:0] iffcq31txctrl0;
wire [15:0] iffcq31txctrl1;
wire [31:0] iffcq31dmonout;
wire [7:0]  iffcq31rxctrl2;
wire [7:0]  iffcq31rxctrl3;
wire [7:0]  iffcq31txctrl2;
wire [1:0]  iffcq31txdeemph;
wire [11:0] iffcq31bufgtdiv;
wire [15:0] iffcq31pinrsrvd;
wire [2:0]  iffcq31loopback;
wire [2:0]  iffcq31rxstatus;
wire [2:0]  iffcq31txmargin;
wire [4:0]  iffcq31txdrvamp;
wire [4:0]  iffcq31txemppos;
wire [4:0]  iffcq31txemppre;
wire [5:0]  iffcq31rxheader;
wire [5:0]  iffcq31txheader;
wire [1:0]  iffcq31refclkpma;
wire [15:0] iffcq31pcsrsvdin;
wire [3:0]  iffcq31rxprbssel;
wire [3:0]  iffcq31txprbssel;
wire [4:0]  iffcq31rxchbondi;
wire [4:0]  iffcq31rxchbondo;
wire [6:0]  iffcq31txempmain;
wire [1:0]  iffcq31rxckcorcnt;
wire [15:0] iffcq31pcsrsvdout;
wire [15:0] iffcq31pinrsrvdas;
wire [6:0]  iffcq31txsequence;
wire [1:0]  iffcq31rxdatavalid;
wire [1:0]  iffcq31rxpowerdown;
wire [1:0]  iffcq31rxresetmode;
wire [1:0]  iffcq31txbufstatus;
wire [1:0]  iffcq31txpowerdown;
wire [1:0]  iffcq31txresetmode;
wire [2:0]  iffcq31rxbufstatus;
wire [3:0]  iffcq31bufgtcemask;
wire [4:0]  iffcq31stepsizeppm;
wire [1:0]  iffcq31rxstartofseq;
wire [3:0]  iffcq31bufgtrstmask;
wire [1:0]  iffcq31rxheadervalid;
wire [2:0]  iffcq31txpmaresetmask;
wire [4:0]  iffcq31rxpcsresetmask;
wire [6:0]  iffcq31rxpmaresetmask;
wire [1:0]  iffcq31rxdapiresetmask;
wire [1:0]  iffcq31txdapiresetmask;
wire [1:0]  iffcq31rxchicoresetmask;
wire [1:0]  iffcq31txchicoresetmask;
wire [7:0]  iffcq31rxethernetstatout;

wire iffcq32enppm;
wire iffcq32perstb;
wire iffcq32bufgtce;
wire iffcq32cdrhold;
wire iffcq32cdrlock;
wire iffcq32dmonclk;
wire iffcq32rxlpmen;
wire iffcq32rxpkdet;
wire iffcq32rxqpien;
wire iffcq32rxslide;
wire iffcq32rxvalid;
wire iffcq32tstclk0;
wire iffcq32tstclk1;
wire iffcq32txswing;
wire iffcq32bufgtrst;
wire iffcq32cdrovren;
wire iffcq32cfokdone;
wire iffcq32iloreset;
wire iffcq32phyready;
wire iffcq32rxlatclk;
wire iffcq32rxusrclk;
wire iffcq32rxusrrdy;
wire iffcq32txcomsas;
wire iffcq32txlatclk;
wire iffcq32txusrclk;
wire iffcq32txusrrdy;
wire iffcq32bsrserial;
wire iffcq32cdrfreqos;
wire iffcq32cdrstepsq;
wire iffcq32cdrstepsx;
wire iffcq32comsasdet;
wire iffcq32gtrxreset;
wire iffcq32gttxreset;
wire iffcq32phystatus;
wire iffcq32rxprbserr;
wire iffcq32rxqpisenn;
wire iffcq32rxqpisenp;
wire iffcq32txcominit;
wire iffcq32txcomwake;
wire iffcq32txdccdone;
wire iffcq32txinhibit;
wire iffcq32txqpisenn;
wire iffcq32txqpisenp;
wire iffcq32aptexthold;
wire iffcq32cdrbmcdreq;
wire iffcq32cdrphreset;
wire iffcq32cdrstepdir;
wire iffcq32cominitdet;
wire iffcq32comwakedet;
wire iffcq32rxcommadet;
wire iffcq32rxelecidle;
wire iffcq32rxoobreset;
wire iffcq32rxpolarity;
wire iffcq32rxsliderdy;
wire iffcq32rxslipdone;
wire iffcq32rxsyncdone;
wire iffcq32txelecidle;
wire iffcq32txpolarity;
wire iffcq32txserpwrdn;
wire iffcq32txsyncdone;
wire iffcq32aptoverwren;
wire iffcq32cdrincpctrl;
wire iffcq32ckpinrsrvd0;
wire iffcq32ckpinrsrvd1;
wire iffcq32cssdstopclk;
wire iffcq32rxcdrphdone;
wire iffcq32rxdapireset;
wire iffcq32rxoutpcsclk;
wire iffcq32rxresetdone;
wire iffcq32rxsyncallin;
wire iffcq32txcomfinish;
wire iffcq32txdapireset;
wire iffcq32txoneszeros;
wire iffcq32txoutpcsclk;
wire iffcq32txqpibiasen;
wire iffcq32txqpiweakpu;
wire iffcq32txresetdone;
wire iffcq32txsyncallin;
wire iffcq32eyescanreset;
wire iffcq32hsdppcsreset;
wire iffcq32iloresetdone;
wire iffcq32iloresetmask;
wire iffcq32rxeqtraining;
wire iffcq32rxphdlyreset;
wire iffcq32rxprbslocked;
wire iffcq32txphdlyreset;
wire iffcq32dmonfiforeset;
wire iffcq32rxbyterealign;
wire iffcq32rxchanbondseq;
wire iffcq32rxchanrealign;
wire iffcq32rxchisaligned;
wire iffcq32rxgearboxslip;
wire iffcq32rxmldchainreq;
wire iffcq32rxtermination;
wire iffcq32txmldchainreq;
wire iffcq32txswingoutlow;
wire iffcq32eyescantrigger;
wire iffcq32resetexception;
wire iffcq32rxmldchaindone;
wire iffcq32rxphasealignpd;
wire iffcq32rxpmaresetdone;
wire iffcq32rxprbscntreset;
wire iffcq32rxprogdivreset;
wire iffcq32tcoclkfsmfrout;
wire iffcq32txchicooutrsvd;
wire iffcq32txmldchaindone;
wire iffcq32txpcsresetmask;
wire iffcq32txphasealignpd;
wire iffcq32txpmaresetdone;
wire iffcq32txprbsforceerr;
wire iffcq32txprogdivreset;
wire iffcq32txswingouthigh;
wire iffcq32rxbyteisaligned;
wire iffcq32rxdapicodereset;
wire iffcq32rxdapiresetdone;
wire iffcq32rxdelayalignerr;
wire iffcq32rxdelayalignreq;
wire iffcq32rxfinealigndone;
wire iffcq32rxphasealignerr;
wire iffcq32rxphasealignreq;
wire iffcq32txdapicodereset;
wire iffcq32txdapiresetdone;
wire iffcq32txdelayalignerr;
wire iffcq32txdelayalignreq;
wire iffcq32txphasealignerr;
wire iffcq32txphasealignreq;
wire iffcq32txtxpicodereset;
wire iffcq32eyescandataerror;
wire iffcq32rxdapicodeovrden;
wire iffcq32rxmlfinealignreq;
wire iffcq32rxphasealigndone;
wire iffcq32txdapicodeovrden;
wire iffcq32txphasealigndone;
wire iffcq32txtxpicodeovrden;
wire iffcq32xpipe5pipelineen;
wire iffcq32rxphasesetinitreq;
wire iffcq32txpausedelayalign;
wire iffcq32txphasesetinitreq;
wire iffcq32rxphasesetinitdone;
wire iffcq32rxphaseshift180req;
wire iffcq32rxprogdivresetdone;
wire iffcq32rxsimplexphystatus;
wire iffcq32txdetectrxloopback;
wire iffcq32txphasesetinitdone;
wire iffcq32txphaseshift180req;
wire iffcq32txprogdivresetdone;
wire iffcq32txsimplexphystatus;
wire iffcq32rxphaseshift180done;
wire iffcq32txphaseshift180done;
wire iffcq32phyesmadaptationsave;
wire iffcq32rxdelayalignprogress;
wire iffcq32txdelayalignprogress;
wire iffcq32rxphasedelayresetdone;
wire iffcq32txphasedelayresetdone;
wire iffcq32txethernetstattxlocalfault;

wire [7:0]  iffcq32rxrate;
wire [7:0]  iffcq32txrate;
wire[127:0] iffcq32rxdata;
wire[127:0] iffcq32txdata;
wire [15:0] iffcq32rxctrl0;
wire [15:0] iffcq32rxctrl1;
wire [15:0] iffcq32txctrl0;
wire [15:0] iffcq32txctrl1;
wire [31:0] iffcq32dmonout;
wire [7:0]  iffcq32rxctrl2;
wire [7:0]  iffcq32rxctrl3;
wire [7:0]  iffcq32txctrl2;
wire [1:0]  iffcq32txdeemph;
wire [11:0] iffcq32bufgtdiv;
wire [15:0] iffcq32pinrsrvd;
wire [2:0]  iffcq32loopback;
wire [2:0]  iffcq32rxstatus;
wire [2:0]  iffcq32txmargin;
wire [4:0]  iffcq32txdrvamp;
wire [4:0]  iffcq32txemppos;
wire [4:0]  iffcq32txemppre;
wire [5:0]  iffcq32rxheader;
wire [5:0]  iffcq32txheader;
wire [1:0]  iffcq32refclkpma;
wire [15:0] iffcq32pcsrsvdin;
wire [3:0]  iffcq32rxprbssel;
wire [3:0]  iffcq32txprbssel;
wire [4:0]  iffcq32rxchbondi;
wire [4:0]  iffcq32rxchbondo;
wire [6:0]  iffcq32txempmain;
wire [1:0]  iffcq32rxckcorcnt;
wire [15:0] iffcq32pcsrsvdout;
wire [15:0] iffcq32pinrsrvdas;
wire [6:0]  iffcq32txsequence;
wire [1:0]  iffcq32rxdatavalid;
wire [1:0]  iffcq32rxpowerdown;
wire [1:0]  iffcq32rxresetmode;
wire [1:0]  iffcq32txbufstatus;
wire [1:0]  iffcq32txpowerdown;
wire [1:0]  iffcq32txresetmode;
wire [2:0]  iffcq32rxbufstatus;
wire [3:0]  iffcq32bufgtcemask;
wire [4:0]  iffcq32stepsizeppm;
wire [1:0]  iffcq32rxstartofseq;
wire [3:0]  iffcq32bufgtrstmask;
wire [1:0]  iffcq32rxheadervalid;
wire [2:0]  iffcq32txpmaresetmask;
wire [4:0]  iffcq32rxpcsresetmask;
wire [6:0]  iffcq32rxpmaresetmask;
wire [1:0]  iffcq32rxdapiresetmask;
wire [1:0]  iffcq32txdapiresetmask;
wire [1:0]  iffcq32rxchicoresetmask;
wire [1:0]  iffcq32txchicoresetmask;
wire [7:0]  iffcq32rxethernetstatout;

wire iffcq33enppm;
wire iffcq33perstb;
wire iffcq33bufgtce;
wire iffcq33cdrhold;
wire iffcq33cdrlock;
wire iffcq33dmonclk;
wire iffcq33rxlpmen;
wire iffcq33rxpkdet;
wire iffcq33rxqpien;
wire iffcq33rxslide;
wire iffcq33rxvalid;
wire iffcq33tstclk0;
wire iffcq33tstclk1;
wire iffcq33txswing;
wire iffcq33bufgtrst;
wire iffcq33cdrovren;
wire iffcq33cfokdone;
wire iffcq33iloreset;
wire iffcq33phyready;
wire iffcq33rxlatclk;
wire iffcq33rxusrclk;
wire iffcq33rxusrrdy;
wire iffcq33txcomsas;
wire iffcq33txlatclk;
wire iffcq33txusrclk;
wire iffcq33txusrrdy;
wire iffcq33bsrserial;
wire iffcq33cdrfreqos;
wire iffcq33cdrstepsq;
wire iffcq33cdrstepsx;
wire iffcq33comsasdet;
wire iffcq33gtrxreset;
wire iffcq33gttxreset;
wire iffcq33phystatus;
wire iffcq33rxprbserr;
wire iffcq33rxqpisenn;
wire iffcq33rxqpisenp;
wire iffcq33txcominit;
wire iffcq33txcomwake;
wire iffcq33txdccdone;
wire iffcq33txinhibit;
wire iffcq33txqpisenn;
wire iffcq33txqpisenp;
wire iffcq33aptexthold;
wire iffcq33cdrbmcdreq;
wire iffcq33cdrphreset;
wire iffcq33cdrstepdir;
wire iffcq33cominitdet;
wire iffcq33comwakedet;
wire iffcq33rxcommadet;
wire iffcq33rxelecidle;
wire iffcq33rxoobreset;
wire iffcq33rxpolarity;
wire iffcq33rxsliderdy;
wire iffcq33rxslipdone;
wire iffcq33rxsyncdone;
wire iffcq33txelecidle;
wire iffcq33txpolarity;
wire iffcq33txserpwrdn;
wire iffcq33txsyncdone;
wire iffcq33aptoverwren;
wire iffcq33cdrincpctrl;
wire iffcq33ckpinrsrvd0;
wire iffcq33ckpinrsrvd1;
wire iffcq33cssdstopclk;
wire iffcq33rxcdrphdone;
wire iffcq33rxdapireset;
wire iffcq33rxoutpcsclk;
wire iffcq33rxresetdone;
wire iffcq33rxsyncallin;
wire iffcq33txcomfinish;
wire iffcq33txdapireset;
wire iffcq33txoneszeros;
wire iffcq33txoutpcsclk;
wire iffcq33txqpibiasen;
wire iffcq33txqpiweakpu;
wire iffcq33txresetdone;
wire iffcq33txsyncallin;
wire iffcq33eyescanreset;
wire iffcq33hsdppcsreset;
wire iffcq33iloresetdone;
wire iffcq33iloresetmask;
wire iffcq33rxeqtraining;
wire iffcq33rxphdlyreset;
wire iffcq33rxprbslocked;
wire iffcq33txphdlyreset;
wire iffcq33dmonfiforeset;
wire iffcq33rxbyterealign;
wire iffcq33rxchanbondseq;
wire iffcq33rxchanrealign;
wire iffcq33rxchisaligned;
wire iffcq33rxgearboxslip;
wire iffcq33rxmldchainreq;
wire iffcq33rxtermination;
wire iffcq33txmldchainreq;
wire iffcq33txswingoutlow;
wire iffcq33eyescantrigger;
wire iffcq33resetexception;
wire iffcq33rxmldchaindone;
wire iffcq33rxphasealignpd;
wire iffcq33rxpmaresetdone;
wire iffcq33rxprbscntreset;
wire iffcq33rxprogdivreset;
wire iffcq33tcoclkfsmfrout;
wire iffcq33txchicooutrsvd;
wire iffcq33txmldchaindone;
wire iffcq33txpcsresetmask;
wire iffcq33txphasealignpd;
wire iffcq33txpmaresetdone;
wire iffcq33txprbsforceerr;
wire iffcq33txprogdivreset;
wire iffcq33txswingouthigh;
wire iffcq33rxbyteisaligned;
wire iffcq33rxdapicodereset;
wire iffcq33rxdapiresetdone;
wire iffcq33rxdelayalignerr;
wire iffcq33rxdelayalignreq;
wire iffcq33rxfinealigndone;
wire iffcq33rxphasealignerr;
wire iffcq33rxphasealignreq;
wire iffcq33txdapicodereset;
wire iffcq33txdapiresetdone;
wire iffcq33txdelayalignerr;
wire iffcq33txdelayalignreq;
wire iffcq33txphasealignerr;
wire iffcq33txphasealignreq;
wire iffcq33txtxpicodereset;
wire iffcq33eyescandataerror;
wire iffcq33rxdapicodeovrden;
wire iffcq33rxmlfinealignreq;
wire iffcq33rxphasealigndone;
wire iffcq33txdapicodeovrden;
wire iffcq33txphasealigndone;
wire iffcq33txtxpicodeovrden;
wire iffcq33xpipe5pipelineen;
wire iffcq33rxphasesetinitreq;
wire iffcq33txpausedelayalign;
wire iffcq33txphasesetinitreq;
wire iffcq33rxphasesetinitdone;
wire iffcq33rxphaseshift180req;
wire iffcq33rxprogdivresetdone;
wire iffcq33rxsimplexphystatus;
wire iffcq33txdetectrxloopback;
wire iffcq33txphasesetinitdone;
wire iffcq33txphaseshift180req;
wire iffcq33txprogdivresetdone;
wire iffcq33txsimplexphystatus;
wire iffcq33rxphaseshift180done;
wire iffcq33txphaseshift180done;
wire iffcq33phyesmadaptationsave;
wire iffcq33rxdelayalignprogress;
wire iffcq33txdelayalignprogress;
wire iffcq33rxphasedelayresetdone;
wire iffcq33txphasedelayresetdone;
wire iffcq33txethernetstattxlocalfault;

wire [7:0]  iffcq33rxrate;
wire [7:0]  iffcq33txrate;
wire[127:0] iffcq33rxdata;
wire[127:0] iffcq33txdata;
wire [15:0] iffcq33rxctrl0;
wire [15:0] iffcq33rxctrl1;
wire [15:0] iffcq33txctrl0;
wire [15:0] iffcq33txctrl1;
wire [31:0] iffcq33dmonout;
wire [7:0]  iffcq33rxctrl2;
wire [7:0]  iffcq33rxctrl3;
wire [7:0]  iffcq33txctrl2;
wire [1:0]  iffcq33txdeemph;
wire [11:0] iffcq33bufgtdiv;
wire [15:0] iffcq33pinrsrvd;
wire [2:0]  iffcq33loopback;
wire [2:0]  iffcq33rxstatus;
wire [2:0]  iffcq33txmargin;
wire [4:0]  iffcq33txdrvamp;
wire [4:0]  iffcq33txemppos;
wire [4:0]  iffcq33txemppre;
wire [5:0]  iffcq33rxheader;
wire [5:0]  iffcq33txheader;
wire [1:0]  iffcq33refclkpma;
wire [15:0] iffcq33pcsrsvdin;
wire [3:0]  iffcq33rxprbssel;
wire [3:0]  iffcq33txprbssel;
wire [4:0]  iffcq33rxchbondi;
wire [4:0]  iffcq33rxchbondo;
wire [6:0]  iffcq33txempmain;
wire [1:0]  iffcq33rxckcorcnt;
wire [15:0] iffcq33pcsrsvdout;
wire [15:0] iffcq33pinrsrvdas;
wire [6:0]  iffcq33txsequence;
wire [1:0]  iffcq33rxdatavalid;
wire [1:0]  iffcq33rxpowerdown;
wire [1:0]  iffcq33rxresetmode;
wire [1:0]  iffcq33txbufstatus;
wire [1:0]  iffcq33txpowerdown;
wire [1:0]  iffcq33txresetmode;
wire [2:0]  iffcq33rxbufstatus;
wire [3:0]  iffcq33bufgtcemask;
wire [4:0]  iffcq33stepsizeppm;
wire [1:0]  iffcq33rxstartofseq;
wire [3:0]  iffcq33bufgtrstmask;
wire [1:0]  iffcq33rxheadervalid;
wire [2:0]  iffcq33txpmaresetmask;
wire [4:0]  iffcq33rxpcsresetmask;
wire [6:0]  iffcq33rxpmaresetmask;
wire [1:0]  iffcq33rxdapiresetmask;
wire [1:0]  iffcq33txdapiresetmask;
wire [1:0]  iffcq33rxchicoresetmask;
wire [1:0]  iffcq33txchicoresetmask;
wire [7:0]  iffcq33rxethernetstatout;

wire iffctrlq0psel;
wire iffctrlq0pready;
wire iffctrlq0pwrite;
wire iffctrlq0apb3clk;
wire iffctrlq0axisclk;
wire iffctrlq0penable;
wire iffctrlq0presetn;
wire iffctrlq0pslverr;
wire iffctrlq0rcalcmp;
wire iffctrlq0rcalenb;
wire iffctrlq0trigin0;
wire iffctrlq0ubmbrst;
wire iffctrlq0bgbypass;
wire iffctrlq0bgpwrdnb;
wire iffctrlq0bgtesten;
wire iffctrlq0trigout0;
wire iffctrlq0ubenable;
wire iffctrlq0ubrxuart;
wire iffctrlq0ubtxuart;
wire iffctrlq0coeregrst;
wire iffctrlq0trigackin0;
wire iffctrlq0ubiolmbrst;
wire iffctrlq0cssdstopclk;
wire iffctrlq0gtpowergood;
wire iffctrlq0m0axistlast;
wire iffctrlq0m1axistlast;
wire iffctrlq0m2axistlast;
wire iffctrlq0rxmarginclk;
wire iffctrlq0s0axistlast;
wire iffctrlq0s1axistlast;
wire iffctrlq0s2axistlast;
wire iffctrlq0trigackout0;
wire iffctrlq0ubinterrupt;
wire iffctrlq0m0axistready;
wire iffctrlq0m0axistvalid;
wire iffctrlq0m1axistready;
wire iffctrlq0m1axistvalid;
wire iffctrlq0m2axistready;
wire iffctrlq0m2axistvalid;
wire iffctrlq0s0axistready;
wire iffctrlq0s0axistvalid;
wire iffctrlq0s1axistready;
wire iffctrlq0s1axistvalid;
wire iffctrlq0s2axistready;
wire iffctrlq0s2axistvalid;
wire iffctrlq0bgrcalovrdenb;
wire iffctrlq0debugtraceclk;
wire iffctrlq0correctableerr;
wire iffctrlq0rxmarginreqack;
wire iffctrlq0rxmarginreqreq;
wire iffctrlq0rxmarginresack;
wire iffctrlq0rxmarginresreq;
wire iffctrlq0debugtracetready;
wire iffctrlq0debugtracetvalid;
wire iffctrlq0uncorrectableerr;
wire iffctrlq0pcielinkreachtarget;

wire [4:0] iffctrlq0rcal;
wire[15:0] iffctrlq0paddr;
wire[31:0] iffctrlq0ubgpi;
wire[31:0] iffctrlq0ubgpo;
wire[11:0] iffctrlq0ubintr;
wire[31:0] iffctrlq0prdata;
wire[31:0] iffctrlq0pwdata;
wire [7:0] iffctrlq0gtrsvdin;
wire [4:0] iffctrlq0bgrcalctl;
wire [7:0] iffctrlq0gtrsvdout;
wire [3:0] iffctrlq0mstrxreset;
wire [3:0] iffctrlq0msttxreset;
wire[31:0] iffctrlq0m0axistdata;
wire[31:0] iffctrlq0m1axistdata;
wire[31:0] iffctrlq0m2axistdata;
wire[31:0] iffctrlq0s0axistdata;
wire[31:0] iffctrlq0s1axistdata;
wire[31:0] iffctrlq0s2axistdata;
wire [3:0] iffctrlq0mstrxresetdone;
wire [3:0] iffctrlq0msttxresetdone;
wire [3:0] iffctrlq0rxmarginreqcmd;
wire [3:0] iffctrlq0rxmarginrescmd;
wire [5:0] iffctrlq0pcieltssmstate;
wire[15:0] iffctrlq0debugtracetdata;
wire [7:0] iffctrlq0rxmarginrespayld;
wire [1:0] iffctrlq0rxmarginreqlanenum;
wire [1:0] iffctrlq0rxmarginreslanenum;
wire [7:0] iffctrlq0rxmarginreqpayload;
wire [7:0] iffctrlq0rxmarginrespayload;

wire iffctrlq1psel;
wire iffctrlq1pready;
wire iffctrlq1pwrite;
wire iffctrlq1apb3clk;
wire iffctrlq1axisclk;
wire iffctrlq1penable;
wire iffctrlq1presetn;
wire iffctrlq1pslverr;
wire iffctrlq1rcalcmp;
wire iffctrlq1rcalenb;
wire iffctrlq1trigin0;
wire iffctrlq1ubmbrst;
wire iffctrlq1bgbypass;
wire iffctrlq1bgpwrdnb;
wire iffctrlq1bgtesten;
wire iffctrlq1trigout0;
wire iffctrlq1ubenable;
wire iffctrlq1ubrxuart;
wire iffctrlq1ubtxuart;
wire iffctrlq1coeregrst;
wire iffctrlq1trigackin0;
wire iffctrlq1ubiolmbrst;
wire iffctrlq1cssdstopclk;
wire iffctrlq1gtpowergood;
wire iffctrlq1m0axistlast;
wire iffctrlq1m1axistlast;
wire iffctrlq1m2axistlast;
wire iffctrlq1rxmarginclk;
wire iffctrlq1s0axistlast;
wire iffctrlq1s1axistlast;
wire iffctrlq1s2axistlast;
wire iffctrlq1trigackout0;
wire iffctrlq1ubinterrupt;
wire iffctrlq1m0axistready;
wire iffctrlq1m0axistvalid;
wire iffctrlq1m1axistready;
wire iffctrlq1m1axistvalid;
wire iffctrlq1m2axistready;
wire iffctrlq1m2axistvalid;
wire iffctrlq1s0axistready;
wire iffctrlq1s0axistvalid;
wire iffctrlq1s1axistready;
wire iffctrlq1s1axistvalid;
wire iffctrlq1s2axistready;
wire iffctrlq1s2axistvalid;
wire iffctrlq1bgrcalovrdenb;
wire iffctrlq1debugtraceclk;
wire iffctrlq1correctableerr;
wire iffctrlq1rxmarginreqack;
wire iffctrlq1rxmarginreqreq;
wire iffctrlq1rxmarginresack;
wire iffctrlq1rxmarginresreq;
wire iffctrlq1debugtracetready;
wire iffctrlq1debugtracetvalid;
wire iffctrlq1uncorrectableerr;
wire iffctrlq1pcielinkreachtarget;

wire [4:0] iffctrlq1rcal;
wire[15:0] iffctrlq1paddr;
wire[31:0] iffctrlq1ubgpi;
wire[31:0] iffctrlq1ubgpo;
wire[11:0] iffctrlq1ubintr;
wire[31:0] iffctrlq1prdata;
wire[31:0] iffctrlq1pwdata;
wire [7:0] iffctrlq1gtrsvdin;
wire [4:0] iffctrlq1bgrcalctl;
wire [7:0] iffctrlq1gtrsvdout;
wire [3:0] iffctrlq1mstrxreset;
wire [3:0] iffctrlq1msttxreset;
wire[31:0] iffctrlq1m0axistdata;
wire[31:0] iffctrlq1m1axistdata;
wire[31:0] iffctrlq1m2axistdata;
wire[31:0] iffctrlq1s0axistdata;
wire[31:0] iffctrlq1s1axistdata;
wire[31:0] iffctrlq1s2axistdata;
wire [3:0] iffctrlq1mstrxresetdone;
wire [3:0] iffctrlq1msttxresetdone;
wire [3:0] iffctrlq1rxmarginreqcmd;
wire [3:0] iffctrlq1rxmarginrescmd;
wire [5:0] iffctrlq1pcieltssmstate;
wire[15:0] iffctrlq1debugtracetdata;
wire [7:0] iffctrlq1rxmarginrespayld;
wire [1:0] iffctrlq1rxmarginreqlanenum;
wire [1:0] iffctrlq1rxmarginreslanenum;
wire [7:0] iffctrlq1rxmarginreqpayload;
wire [7:0] iffctrlq1rxmarginrespayload;

wire iffctrlq2psel;
wire iffctrlq2pready;
wire iffctrlq2pwrite;
wire iffctrlq2apb3clk;
wire iffctrlq2axisclk;
wire iffctrlq2penable;
wire iffctrlq2presetn;
wire iffctrlq2pslverr;
wire iffctrlq2rcalcmp;
wire iffctrlq2rcalenb;
wire iffctrlq2trigin0;
wire iffctrlq2ubmbrst;
wire iffctrlq2bgbypass;
wire iffctrlq2bgpwrdnb;
wire iffctrlq2bgtesten;
wire iffctrlq2trigout0;
wire iffctrlq2ubenable;
wire iffctrlq2ubrxuart;
wire iffctrlq2ubtxuart;
wire iffctrlq2coeregrst;
wire iffctrlq2trigackin0;
wire iffctrlq2ubiolmbrst;
wire iffctrlq2cssdstopclk;
wire iffctrlq2gtpowergood;
wire iffctrlq2m0axistlast;
wire iffctrlq2m1axistlast;
wire iffctrlq2m2axistlast;
wire iffctrlq2rxmarginclk;
wire iffctrlq2s0axistlast;
wire iffctrlq2s1axistlast;
wire iffctrlq2s2axistlast;
wire iffctrlq2trigackout0;
wire iffctrlq2ubinterrupt;
wire iffctrlq2m0axistready;
wire iffctrlq2m0axistvalid;
wire iffctrlq2m1axistready;
wire iffctrlq2m1axistvalid;
wire iffctrlq2m2axistready;
wire iffctrlq2m2axistvalid;
wire iffctrlq2s0axistready;
wire iffctrlq2s0axistvalid;
wire iffctrlq2s1axistready;
wire iffctrlq2s1axistvalid;
wire iffctrlq2s2axistready;
wire iffctrlq2s2axistvalid;
wire iffctrlq2bgrcalovrdenb;
wire iffctrlq2debugtraceclk;
wire iffctrlq2correctableerr;
wire iffctrlq2rxmarginreqack;
wire iffctrlq2rxmarginreqreq;
wire iffctrlq2rxmarginresack;
wire iffctrlq2rxmarginresreq;
wire iffctrlq2debugtracetready;
wire iffctrlq2debugtracetvalid;
wire iffctrlq2uncorrectableerr;
wire iffctrlq2pcielinkreachtarget;

wire [4:0] iffctrlq2rcal;
wire[15:0] iffctrlq2paddr;
wire[31:0] iffctrlq2ubgpi;
wire[31:0] iffctrlq2ubgpo;
wire[11:0] iffctrlq2ubintr;
wire[31:0] iffctrlq2prdata;
wire[31:0] iffctrlq2pwdata;
wire [7:0] iffctrlq2gtrsvdin;
wire [4:0] iffctrlq2bgrcalctl;
wire [7:0] iffctrlq2gtrsvdout;
wire [3:0] iffctrlq2mstrxreset;
wire [3:0] iffctrlq2msttxreset;
wire[31:0] iffctrlq2m0axistdata;
wire[31:0] iffctrlq2m1axistdata;
wire[31:0] iffctrlq2m2axistdata;
wire[31:0] iffctrlq2s0axistdata;
wire[31:0] iffctrlq2s1axistdata;
wire[31:0] iffctrlq2s2axistdata;
wire [3:0] iffctrlq2mstrxresetdone;
wire [3:0] iffctrlq2msttxresetdone;
wire [3:0] iffctrlq2rxmarginreqcmd;
wire [3:0] iffctrlq2rxmarginrescmd;
wire [5:0] iffctrlq2pcieltssmstate;
wire[15:0] iffctrlq2debugtracetdata;
wire [7:0] iffctrlq2rxmarginrespayld;
wire [1:0] iffctrlq2rxmarginreqlanenum;
wire [1:0] iffctrlq2rxmarginreslanenum;
wire [7:0] iffctrlq2rxmarginreqpayload;
wire [7:0] iffctrlq2rxmarginrespayload;

wire iffctrlq3psel;
wire iffctrlq3pready;
wire iffctrlq3pwrite;
wire iffctrlq3apb3clk;
wire iffctrlq3axisclk;
wire iffctrlq3penable;
wire iffctrlq3presetn;
wire iffctrlq3pslverr;
wire iffctrlq3rcalcmp;
wire iffctrlq3rcalenb;
wire iffctrlq3trigin0;
wire iffctrlq3ubmbrst;
wire iffctrlq3bgbypass;
wire iffctrlq3bgpwrdnb;
wire iffctrlq3bgtesten;
wire iffctrlq3trigout0;
wire iffctrlq3ubenable;
wire iffctrlq3ubrxuart;
wire iffctrlq3ubtxuart;
wire iffctrlq3coeregrst;
wire iffctrlq3trigackin0;
wire iffctrlq3ubiolmbrst;
wire iffctrlq3cssdstopclk;
wire iffctrlq3gtpowergood;
wire iffctrlq3m0axistlast;
wire iffctrlq3m1axistlast;
wire iffctrlq3m2axistlast;
wire iffctrlq3rxmarginclk;
wire iffctrlq3s0axistlast;
wire iffctrlq3s1axistlast;
wire iffctrlq3s2axistlast;
wire iffctrlq3trigackout0;
wire iffctrlq3ubinterrupt;
wire iffctrlq3m0axistready;
wire iffctrlq3m0axistvalid;
wire iffctrlq3m1axistready;
wire iffctrlq3m1axistvalid;
wire iffctrlq3m2axistready;
wire iffctrlq3m2axistvalid;
wire iffctrlq3s0axistready;
wire iffctrlq3s0axistvalid;
wire iffctrlq3s1axistready;
wire iffctrlq3s1axistvalid;
wire iffctrlq3s2axistready;
wire iffctrlq3s2axistvalid;
wire iffctrlq3bgrcalovrdenb;
wire iffctrlq3debugtraceclk;
wire iffctrlq3correctableerr;
wire iffctrlq3rxmarginreqack;
wire iffctrlq3rxmarginreqreq;
wire iffctrlq3rxmarginresack;
wire iffctrlq3rxmarginresreq;
wire iffctrlq3debugtracetready;
wire iffctrlq3debugtracetvalid;
wire iffctrlq3uncorrectableerr;
wire iffctrlq3pcielinkreachtarget;

wire [4:0] iffctrlq3rcal;
wire[15:0] iffctrlq3paddr;
wire[31:0] iffctrlq3ubgpi;
wire[31:0] iffctrlq3ubgpo;
wire[11:0] iffctrlq3ubintr;
wire[31:0] iffctrlq3prdata;
wire[31:0] iffctrlq3pwdata;
wire [7:0] iffctrlq3gtrsvdin;
wire [4:0] iffctrlq3bgrcalctl;
wire [7:0] iffctrlq3gtrsvdout;
wire [3:0] iffctrlq3mstrxreset;
wire [3:0] iffctrlq3msttxreset;
wire[31:0] iffctrlq3m0axistdata;
wire[31:0] iffctrlq3m1axistdata;
wire[31:0] iffctrlq3m2axistdata;
wire[31:0] iffctrlq3s0axistdata;
wire[31:0] iffctrlq3s1axistdata;
wire[31:0] iffctrlq3s2axistdata;
wire [3:0] iffctrlq3mstrxresetdone;
wire [3:0] iffctrlq3msttxresetdone;
wire [3:0] iffctrlq3rxmarginreqcmd;
wire [3:0] iffctrlq3rxmarginrescmd;
wire [5:0] iffctrlq3pcieltssmstate;
wire[15:0] iffctrlq3debugtracetdata;
wire [7:0] iffctrlq3rxmarginrespayld;
wire [1:0] iffctrlq3rxmarginreqlanenum;
wire [1:0] iffctrlq3rxmarginreslanenum;
wire [7:0] iffctrlq3rxmarginreqpayload;
wire [7:0] iffctrlq3rxmarginrespayload;

wire iffhsq00rpllpwrdn;
wire iffhsq00rpllreset;
wire iffhsq00lcpllpwrdn;
wire iffhsq00lcpllreset;
wire iffhsq00rpllfbloss;
wire iffhsq00corerefclk0;
wire iffhsq00corerefclk1;
wire iffhsq00lcpllfbloss;
wire iffhsq00rpllrefloss;
wire iffhsq00lcpllrefloss;
wire iffhsq00rpllfreqlock;
wire iffhsq00rxrecclkout0;
wire iffhsq00rxrecclkout1;
wire iffhsq00lcpllfreqlock;
wire iffhsq00rpllsdmtoggle;
wire iffhsq00lcpllsdmtoggle;
wire iffhsq00mgtrpllrefclkfa;
wire iffhsq00mgtlcpllrefclkfa;
wire iffhsq00rpllresetbypassmode;
wire iffhsq00lcpllresetbypassmode;

wire [7:0] iffhsq00rpllfbdiv;
wire [7:0] iffhsq00lcpllfbdiv;
wire[25:0] iffhsq00rpllsdmdata;
wire[25:0] iffhsq00lcpllsdmdata;
wire [1:0] iffhsq00rpllresetmask;
wire [2:0] iffhsq00rpllrefseldyn;
wire [1:0] iffhsq00lcpllresetmask;
wire [2:0] iffhsq00lcpllrefseldyn;

wire iffhsq01rpllpwrdn;
wire iffhsq01rpllreset;
wire iffhsq01lcpllpwrdn;
wire iffhsq01lcpllreset;
wire iffhsq01rpllfbloss;
wire iffhsq01corerefclk0;
wire iffhsq01corerefclk1;
wire iffhsq01lcpllfbloss;
wire iffhsq01rpllrefloss;
wire iffhsq01lcpllrefloss;
wire iffhsq01rxrecclkout0;
wire iffhsq01rxrecclkout1;
wire iffhsq01rpllfreqlock;
wire iffhsq01lcpllfreqlock;
wire iffhsq01rpllsdmtoggle;
wire iffhsq01lcpllsdmtoggle;
wire iffhsq01mgtrpllrefclkfa;
wire iffhsq01mgtlcpllrefclkfa;
wire iffhsq01rpllresetbypassmode;
wire iffhsq01lcpllresetbypassmode;

wire [7:0] iffhsq01rpllfbdiv;
wire [7:0] iffhsq01lcpllfbdiv;
wire[25:0] iffhsq01rpllsdmdata;
wire[25:0] iffhsq01lcpllsdmdata;
wire [1:0] iffhsq01rpllresetmask;
wire [2:0] iffhsq01rpllrefseldyn;
wire [1:0] iffhsq01lcpllresetmask;
wire [2:0] iffhsq01lcpllrefseldyn;

wire iffhsq10rpllpwrdn;
wire iffhsq10rpllreset;
wire iffhsq10lcpllpwrdn;
wire iffhsq10lcpllreset;
wire iffhsq10rpllfbloss;
wire iffhsq10corerefclk0;
wire iffhsq10corerefclk1;
wire iffhsq10lcpllfbloss;
wire iffhsq10rpllrefloss;
wire iffhsq10lcpllrefloss;
wire iffhsq10rxrecclkout0;
wire iffhsq10rxrecclkout1;
wire iffhsq10rpllfreqlock;
wire iffhsq10lcpllfreqlock;
wire iffhsq10rpllsdmtoggle;
wire iffhsq10lcpllsdmtoggle;
wire iffhsq10mgtrpllrefclkfa;
wire iffhsq10mgtlcpllrefclkfa;
wire iffhsq10rpllresetbypassmode;
wire iffhsq10lcpllresetbypassmode;

wire [7:0] iffhsq10rpllfbdiv;
wire [7:0] iffhsq10lcpllfbdiv;
wire[25:0] iffhsq10rpllsdmdata;
wire[25:0] iffhsq10lcpllsdmdata;
wire [1:0] iffhsq10rpllresetmask;
wire [2:0] iffhsq10rpllrefseldyn;
wire [1:0] iffhsq10lcpllresetmask;
wire [2:0] iffhsq10lcpllrefseldyn;

wire iffhsq11rpllpwrdn;
wire iffhsq11rpllreset;
wire iffhsq11lcpllpwrdn;
wire iffhsq11lcpllreset;
wire iffhsq11rpllfbloss;
wire iffhsq11corerefclk0;
wire iffhsq11corerefclk1;
wire iffhsq11lcpllfbloss;
wire iffhsq11rpllrefloss;
wire iffhsq11lcpllrefloss;
wire iffhsq11rpllfreqlock;
wire iffhsq11rxrecclkout0;
wire iffhsq11rxrecclkout1;
wire iffhsq11lcpllfreqlock;
wire iffhsq11rpllsdmtoggle;
wire iffhsq11lcpllsdmtoggle;
wire iffhsq11mgtrpllrefclkfa;
wire iffhsq11mgtlcpllrefclkfa;
wire iffhsq11rpllresetbypassmode;
wire iffhsq11lcpllresetbypassmode;

wire [7:0] iffhsq11rpllfbdiv;
wire [7:0] iffhsq11lcpllfbdiv;
wire[25:0] iffhsq11rpllsdmdata;
wire[25:0] iffhsq11lcpllsdmdata;
wire [1:0] iffhsq11rpllresetmask;
wire [2:0] iffhsq11rpllrefseldyn;
wire [1:0] iffhsq11lcpllresetmask;
wire [2:0] iffhsq11lcpllrefseldyn;

wire iffhsq20rpllpwrdn;
wire iffhsq20rpllreset;
wire iffhsq20lcpllpwrdn;
wire iffhsq20lcpllreset;
wire iffhsq20rpllfbloss;
wire iffhsq20corerefclk0;
wire iffhsq20corerefclk1;
wire iffhsq20lcpllfbloss;
wire iffhsq20rpllrefloss;
wire iffhsq20lcpllrefloss;
wire iffhsq20rpllfreqlock;
wire iffhsq20rxrecclkout0;
wire iffhsq20rxrecclkout1;
wire iffhsq20lcpllfreqlock;
wire iffhsq20rpllsdmtoggle;
wire iffhsq20lcpllsdmtoggle;
wire iffhsq20mgtrpllrefclkfa;
wire iffhsq20mgtlcpllrefclkfa;
wire iffhsq20rpllresetbypassmode;
wire iffhsq20lcpllresetbypassmode;

wire [7:0] iffhsq20rpllfbdiv;
wire [7:0] iffhsq20lcpllfbdiv;
wire[25:0] iffhsq20rpllsdmdata;
wire[25:0] iffhsq20lcpllsdmdata;
wire [1:0] iffhsq20rpllresetmask;
wire [2:0] iffhsq20rpllrefseldyn;
wire [1:0] iffhsq20lcpllresetmask;
wire [2:0] iffhsq20lcpllrefseldyn;

wire iffhsq21rpllpwrdn;
wire iffhsq21rpllreset;
wire iffhsq21lcpllpwrdn;
wire iffhsq21lcpllreset;
wire iffhsq21rpllfbloss;
wire iffhsq21corerefclk0;
wire iffhsq21corerefclk1;
wire iffhsq21lcpllfbloss;
wire iffhsq21rpllrefloss;
wire iffhsq21lcpllrefloss;
wire iffhsq21rpllfreqlock;
wire iffhsq21rxrecclkout0;
wire iffhsq21rxrecclkout1;
wire iffhsq21lcpllfreqlock;
wire iffhsq21rpllsdmtoggle;
wire iffhsq21lcpllsdmtoggle;
wire iffhsq21mgtrpllrefclkfa;
wire iffhsq21mgtlcpllrefclkfa;
wire iffhsq21rpllresetbypassmode;
wire iffhsq21lcpllresetbypassmode;

wire [7:0] iffhsq21rpllfbdiv;
wire [7:0] iffhsq21lcpllfbdiv;
wire[25:0] iffhsq21rpllsdmdata;
wire[25:0] iffhsq21lcpllsdmdata;
wire [1:0] iffhsq21rpllresetmask;
wire [2:0] iffhsq21rpllrefseldyn;
wire [1:0] iffhsq21lcpllresetmask;
wire [2:0] iffhsq21lcpllrefseldyn;

wire iffhsq30rpllpwrdn;
wire iffhsq30rpllreset;
wire iffhsq30lcpllpwrdn;
wire iffhsq30lcpllreset;
wire iffhsq30rpllfbloss;
wire iffhsq30corerefclk0;
wire iffhsq30corerefclk1;
wire iffhsq30lcpllfbloss;
wire iffhsq30rpllrefloss;
wire iffhsq30lcpllrefloss;
wire iffhsq30rpllfreqlock;
wire iffhsq30rxrecclkout0;
wire iffhsq30rxrecclkout1;
wire iffhsq30lcpllfreqlock;
wire iffhsq30rpllsdmtoggle;
wire iffhsq30lcpllsdmtoggle;
wire iffhsq30mgtrpllrefclkfa;
wire iffhsq30mgtlcpllrefclkfa;
wire iffhsq30rpllresetbypassmode;
wire iffhsq30lcpllresetbypassmode;

wire [7:0] iffhsq30rpllfbdiv;
wire [7:0] iffhsq30lcpllfbdiv;
wire[25:0] iffhsq30rpllsdmdata;
wire[25:0] iffhsq30lcpllsdmdata;
wire [1:0] iffhsq30rpllresetmask;
wire [2:0] iffhsq30rpllrefseldyn;
wire [1:0] iffhsq30lcpllresetmask;
wire [2:0] iffhsq30lcpllrefseldyn;

wire iffhsq31rpllpwrdn;
wire iffhsq31rpllreset;
wire iffhsq31lcpllpwrdn;
wire iffhsq31lcpllreset;
wire iffhsq31rpllfbloss;
wire iffhsq31corerefclk0;
wire iffhsq31corerefclk1;
wire iffhsq31lcpllfbloss;
wire iffhsq31rpllrefloss;
wire iffhsq31lcpllrefloss;
wire iffhsq31rpllfreqlock;
wire iffhsq31rxrecclkout0;
wire iffhsq31rxrecclkout1;
wire iffhsq31lcpllfreqlock;
wire iffhsq31rpllsdmtoggle;
wire iffhsq31lcpllsdmtoggle;
wire iffhsq31mgtrpllrefclkfa;
wire iffhsq31mgtlcpllrefclkfa;
wire iffhsq31rpllresetbypassmode;
wire iffhsq31lcpllresetbypassmode;

wire [7:0] iffhsq31rpllfbdiv;
wire [7:0] iffhsq31lcpllfbdiv;
wire[25:0] iffhsq31rpllsdmdata;
wire[25:0] iffhsq31lcpllsdmdata;
wire [1:0] iffhsq31rpllresetmask;
wire [2:0] iffhsq31rpllrefseldyn;
wire [1:0] iffhsq31lcpllresetmask;
wire [2:0] iffhsq31lcpllrefseldyn;

wire iffrckq00refclkpd;
wire iffrckq01refclkpd;
wire iffrckq10refclkpd;
wire iffrckq11refclkpd;
wire iffrckq20refclkpd;
wire iffrckq21refclkpd;
wire iffrckq30refclkpd;
wire iffrckq31refclkpd;
wire iffrckq00hrowtestck;
wire iffrckq01hrowtestck;
wire iffrckq10hrowtestck;
wire iffrckq11hrowtestck;
wire iffrckq20hrowtestck;
wire iffrckq21hrowtestck;
wire iffrckq30hrowtestck;
wire iffrckq31hrowtestck;

wire ifplcpm5p0chimsactive;
wire ifplcpm5p0chireqflitv;
wire ifplcpm5p0chireqlcrdv;
wire ifplcpm5p0chisnpflitv;
wire ifplcpm5p0chisnplcrdv;
wire ifplcpm5p0chissactive;
wire ifplcpm5p0chisyscoack;
wire ifplcpm5p0chisyscoreq;
wire ifplcpm5p0chicrspflitv;
wire ifplcpm5p0chicrsplcrdv;
wire ifplcpm5p0chirdatflitv;
wire ifplcpm5p0chirdatlcrdv;
wire ifplcpm5p0chisrspflitv;
wire ifplcpm5p0chisrsplcrdv;
wire ifplcpm5p0chiwdatflitv;
wire ifplcpm5p0chiwdatlcrdv;
wire ifplcpm5p0chireqflitpend;
wire ifplcpm5p0chisnpflitpend;
wire ifplcpm5p0chicrspflitpend;
wire ifplcpm5p0chirdatflitpend;
wire ifplcpm5p0chisrspflitpend;
wire ifplcpm5p0chiwdatflitpend;
wire ifplcpm5p0chimlinkactiveack;
wire ifplcpm5p0chimlinkactivereq;
wire ifplcpm5p0chislinkactiveack;
wire ifplcpm5p0chislinkactivereq;

wire [87:0] ifplcpm5p0chisnpflit;
wire[120:0] ifplcpm5p0chireqflit;
wire [50:0] ifplcpm5p0chicrspflit;
wire [50:0] ifplcpm5p0chisrspflit;
wire[704:0] ifplcpm5p0chirdatflit;
wire[704:0] ifplcpm5p0chiwdatflit;

wire ifplcpm5p1chimsactive;
wire ifplcpm5p1chireqflitv;
wire ifplcpm5p1chireqlcrdv;
wire ifplcpm5p1chisnpflitv;
wire ifplcpm5p1chisnplcrdv;
wire ifplcpm5p1chissactive;
wire ifplcpm5p1chisyscoack;
wire ifplcpm5p1chisyscoreq;
wire ifplcpm5p1chicrspflitv;
wire ifplcpm5p1chicrsplcrdv;
wire ifplcpm5p1chirdatflitv;
wire ifplcpm5p1chirdatlcrdv;
wire ifplcpm5p1chisrspflitv;
wire ifplcpm5p1chisrsplcrdv;
wire ifplcpm5p1chiwdatflitv;
wire ifplcpm5p1chiwdatlcrdv;
wire ifplcpm5p1chireqflitpend;
wire ifplcpm5p1chisnpflitpend;
wire ifplcpm5p1chicrspflitpend;
wire ifplcpm5p1chirdatflitpend;
wire ifplcpm5p1chisrspflitpend;
wire ifplcpm5p1chiwdatflitpend;
wire ifplcpm5p1chimlinkactiveack;
wire ifplcpm5p1chimlinkactivereq;
wire ifplcpm5p1chislinkactiveack;
wire ifplcpm5p1chislinkactivereq;

wire [87:0] ifplcpm5p1chisnpflit;
wire[120:0] ifplcpm5p1chireqflit;
wire [50:0] ifplcpm5p1chicrspflit;
wire [50:0] ifplcpm5p1chisrspflit;
wire[704:0] ifplcpm5p1chirdatflit;
wire[704:0] ifplcpm5p1chiwdatflit;

wire ifpscpmchannel0xpiperxvalid;
wire ifpscpmchannel0xpipephystatus;
wire ifpscpmchannel0xpiperxelecidle;
wire ifpscpmchannel0xpiperxdatavalid;
wire ifpscpmchannel0xpiperxstartblock;
wire[31:0] ifpscpmchannel0xpiperxdata;
wire [2:0] ifpscpmchannel0xpiperxstatus;
wire [1:0] ifpscpmchannel0xpiperxcharisk;
wire [1:0] ifpscpmchannel0xpiperxsyncheader;

wire ifpscpmchannel1xpiperxvalid;
wire ifpscpmchannel1xpipephystatus;
wire ifpscpmchannel1xpiperxelecidle;
wire ifpscpmchannel1xpiperxdatavalid;
wire ifpscpmchannel1xpiperxstartblock;
wire[31:0] ifpscpmchannel1xpiperxdata;
wire [2:0] ifpscpmchannel1xpiperxstatus;
wire [1:0] ifpscpmchannel1xpiperxcharisk;
wire [1:0] ifpscpmchannel1xpiperxsyncheader;

wire ifpscpmchannel2xpiperxvalid;
wire ifpscpmchannel2xpipephystatus;
wire ifpscpmchannel2xpiperxelecidle;
wire ifpscpmchannel2xpiperxdatavalid;
wire ifpscpmchannel2xpiperxstartblock;
wire[31:0] ifpscpmchannel2xpiperxdata;
wire [2:0] ifpscpmchannel2xpiperxstatus;
wire [1:0] ifpscpmchannel2xpiperxcharisk;
wire [1:0] ifpscpmchannel2xpiperxsyncheader;

wire ifpscpmchannel3xpiperxvalid;
wire ifpscpmchannel3xpipephystatus;
wire ifpscpmchannel3xpiperxelecidle;
wire ifpscpmchannel3xpiperxdatavalid;
wire ifpscpmchannel3xpiperxstartblock;
wire[31:0] ifpscpmchannel3xpiperxdata;
wire [2:0] ifpscpmchannel3xpiperxstatus;
wire [1:0] ifpscpmchannel3xpiperxcharisk;
wire [1:0] ifpscpmchannel3xpiperxsyncheader;

wire ifpscpmchannel4xpiperxvalid;
wire ifpscpmchannel4xpipephystatus;
wire ifpscpmchannel4xpiperxelecidle;
wire ifpscpmchannel4xpiperxdatavalid;
wire ifpscpmchannel4xpiperxstartblock;
wire[31:0] ifpscpmchannel4xpiperxdata;
wire [2:0] ifpscpmchannel4xpiperxstatus;
wire [1:0] ifpscpmchannel4xpiperxcharisk;
wire [1:0] ifpscpmchannel4xpiperxsyncheader;

wire ifpscpmchannel5xpiperxvalid;
wire ifpscpmchannel5xpipephystatus;
wire ifpscpmchannel5xpiperxelecidle;
wire ifpscpmchannel5xpiperxdatavalid;
wire ifpscpmchannel5xpiperxstartblock;
wire[31:0] ifpscpmchannel5xpiperxdata;
wire [2:0] ifpscpmchannel5xpiperxstatus;
wire [1:0] ifpscpmchannel5xpiperxcharisk;
wire [1:0] ifpscpmchannel5xpiperxsyncheader;

wire ifpscpmchannel6xpiperxvalid;
wire ifpscpmchannel6xpipephystatus;
wire ifpscpmchannel6xpiperxelecidle;
wire ifpscpmchannel6xpiperxdatavalid;
wire ifpscpmchannel6xpiperxstartblock;
wire[31:0] ifpscpmchannel6xpiperxdata;
wire [2:0] ifpscpmchannel6xpiperxstatus;
wire [1:0] ifpscpmchannel6xpiperxcharisk;
wire [1:0] ifpscpmchannel6xpiperxsyncheader;

wire ifpscpmchannel7xpiperxvalid;
wire ifpscpmchannel7xpipephystatus;
wire ifpscpmchannel7xpiperxelecidle;
wire ifpscpmchannel7xpiperxdatavalid;
wire ifpscpmchannel7xpiperxstartblock;
wire[31:0] ifpscpmchannel7xpiperxdata;
wire [2:0] ifpscpmchannel7xpiperxstatus;
wire [1:0] ifpscpmchannel7xpiperxcharisk;
wire [1:0] ifpscpmchannel7xpiperxsyncheader;

wire ifpscpmchannel8xpiperxvalid;
wire ifpscpmchannel8xpipephystatus;
wire ifpscpmchannel8xpiperxelecidle;
wire ifpscpmchannel8xpiperxdatavalid;
wire ifpscpmchannel8xpiperxstartblock;
wire[31:0] ifpscpmchannel8xpiperxdata;
wire [2:0] ifpscpmchannel8xpiperxstatus;
wire [1:0] ifpscpmchannel8xpiperxcharisk;
wire [1:0] ifpscpmchannel8xpiperxsyncheader;

wire ifpscpmchannel9xpiperxvalid;
wire ifpscpmchannel9xpipephystatus;
wire ifpscpmchannel9xpiperxelecidle;
wire ifpscpmchannel9xpiperxdatavalid;
wire ifpscpmchannel9xpiperxstartblock;
wire[31:0] ifpscpmchannel9xpiperxdata;
wire [2:0] ifpscpmchannel9xpiperxstatus;
wire [1:0] ifpscpmchannel9xpiperxcharisk;
wire [1:0] ifpscpmchannel9xpiperxsyncheader;

wire ifpscpmchannel10xpiperxvalid;
wire ifpscpmchannel10xpipephystatus;
wire ifpscpmchannel10xpiperxelecidle;
wire ifpscpmchannel10xpiperxdatavalid;
wire ifpscpmchannel10xpiperxstartblock;
wire[31:0] ifpscpmchannel10xpiperxdata;
wire [2:0] ifpscpmchannel10xpiperxstatus;
wire [1:0] ifpscpmchannel10xpiperxcharisk;
wire [1:0] ifpscpmchannel10xpiperxsyncheader;

wire ifpscpmchannel11xpiperxvalid;
wire ifpscpmchannel11xpipephystatus;
wire ifpscpmchannel11xpiperxelecidle;
wire ifpscpmchannel11xpiperxdatavalid;
wire ifpscpmchannel11xpiperxstartblock;
wire[31:0] ifpscpmchannel11xpiperxdata;
wire [2:0] ifpscpmchannel11xpiperxstatus;
wire [1:0] ifpscpmchannel11xpiperxcharisk;
wire [1:0] ifpscpmchannel11xpiperxsyncheader;

wire ifpscpmchannel12xpiperxvalid;
wire ifpscpmchannel12xpipephystatus;
wire ifpscpmchannel12xpiperxelecidle;
wire ifpscpmchannel12xpiperxdatavalid;
wire ifpscpmchannel12xpiperxstartblock;
wire[31:0] ifpscpmchannel12xpiperxdata;
wire [2:0] ifpscpmchannel12xpiperxstatus;
wire [1:0] ifpscpmchannel12xpiperxcharisk;
wire [1:0] ifpscpmchannel12xpiperxsyncheader;

wire ifpscpmchannel13xpiperxvalid;
wire ifpscpmchannel13xpipephystatus;
wire ifpscpmchannel13xpiperxelecidle;
wire ifpscpmchannel13xpiperxdatavalid;
wire ifpscpmchannel13xpiperxstartblock;
wire[31:0] ifpscpmchannel13xpiperxdata;
wire [2:0] ifpscpmchannel13xpiperxstatus;
wire [1:0] ifpscpmchannel13xpiperxcharisk;
wire [1:0] ifpscpmchannel13xpiperxsyncheader;

wire ifpscpmchannel14xpiperxvalid;
wire ifpscpmchannel14xpipephystatus;
wire ifpscpmchannel14xpiperxelecidle;
wire ifpscpmchannel14xpiperxdatavalid;
wire ifpscpmchannel14xpiperxstartblock;
wire[31:0] ifpscpmchannel14xpiperxdata;
wire [2:0] ifpscpmchannel14xpiperxstatus;
wire [1:0] ifpscpmchannel14xpiperxcharisk;
wire [1:0] ifpscpmchannel14xpiperxsyncheader;

wire ifpscpmchannel15xpiperxvalid;
wire ifpscpmchannel15xpipephystatus;
wire ifpscpmchannel15xpiperxelecidle;
wire ifpscpmchannel15xpiperxdatavalid;
wire ifpscpmchannel15xpiperxstartblock;
wire[31:0] ifpscpmchannel15xpiperxdata;
wire [2:0] ifpscpmchannel15xpiperxstatus;
wire [1:0] ifpscpmchannel15xpiperxcharisk;
wire [1:0] ifpscpmchannel15xpiperxsyncheader;

wire ifpscpmhsdpchannel0xpiperxdatavalid;
wire ifpscpmhsdpchannel0xpiperxresetdone;
wire ifpscpmhsdpchannel0xpipetxresetdone;
wire ifpscpmhsdpchannel1xpiperxdatavalid;
wire ifpscpmhsdpchannel1xpiperxresetdone;
wire ifpscpmhsdpchannel1xpipetxresetdone;
wire ifpscpmhsdpchannel2xpiperxdatavalid;
wire ifpscpmhsdpchannel2xpiperxresetdone;
wire ifpscpmhsdpchannel2xpipetxresetdone;
wire ifpscpmhsdpchannel0xpiperxheadervalid;
wire ifpscpmhsdpchannel1xpiperxheadervalid;
wire ifpscpmhsdpchannel2xpiperxheadervalid;
wire [1:0] ifpscpmhsdpchannel0xpiperxheader;
wire [1:0] ifpscpmhsdpchannel1xpiperxheader;
wire [1:0] ifpscpmhsdpchannel2xpiperxheader;

wire ifpscpmhsdplinkxpipegtrxoutclk;

wire ifpscpmlink0xpipebufgtce;
wire ifpscpmlink0xpipebufgtrst;
wire ifpscpmlink0xpipegtoutclk;
wire ifpscpmlink0xpipephyready;
wire ifpscpmlink1xpipebufgtce;
wire ifpscpmlink1xpipebufgtrst;
wire ifpscpmlink1xpipegtoutclk;
wire ifpscpmlink1xpipephyready;
wire[11:0] ifpscpmlink0xpipebufgtdiv;
wire[11:0] ifpscpmlink1xpipebufgtdiv;
wire [3:0] ifpscpmlink0xpipebufgtcemask;
wire [3:0] ifpscpmlink1xpipebufgtcemask;
wire [3:0] ifpscpmlink0xpipebufgtrstmask;
wire [3:0] ifpscpmlink1xpipebufgtrstmask;

wire ifpscpmintquadxpipephyreadytobot;

wire ifpscpmpcsrpsrincal;
wire ifpscpmpcsrpsrbisrerr;
wire ifpscpmpcsrpsrcaldone;
wire ifpscpmpcsrpsrbisrdone;
wire ifpscpmpcsrpsrcalerror;
wire ifpscpmpcsrpsrmemclrdone;
wire ifpscpmpcsrpsrmemclrpass;
wire ifpscpmpcsrpsrscanclrdone;
wire ifpscpmpcsrpsrscanclrpass;

wire ifpscpmquad0xpiperxmarginreqack;
wire ifpscpmquad0xpiperxmarginreqreq;
wire ifpscpmquad0xpiperxmarginresack;
wire ifpscpmquad0xpiperxmarginresreq;
wire ifpscpmquad1xpiperxmarginreqack;
wire ifpscpmquad1xpiperxmarginreqreq;
wire ifpscpmquad1xpiperxmarginresack;
wire ifpscpmquad1xpiperxmarginresreq;
wire ifpscpmquad2xpiperxmarginreqack;
wire ifpscpmquad2xpiperxmarginreqreq;
wire ifpscpmquad2xpiperxmarginresack;
wire ifpscpmquad2xpiperxmarginresreq;
wire ifpscpmquad3xpiperxmarginreqack;
wire ifpscpmquad3xpiperxmarginreqreq;
wire ifpscpmquad3xpiperxmarginresack;
wire ifpscpmquad3xpiperxmarginresreq;

wire [3:0] ifpscpmquad0xpiperxmarginreqcmd;
wire [3:0] ifpscpmquad0xpiperxmarginrescmd;
wire [3:0] ifpscpmquad1xpiperxmarginreqcmd;
wire [3:0] ifpscpmquad1xpiperxmarginrescmd;
wire [3:0] ifpscpmquad2xpiperxmarginreqcmd;
wire [3:0] ifpscpmquad2xpiperxmarginrescmd;
wire [3:0] ifpscpmquad3xpiperxmarginreqcmd;
wire [3:0] ifpscpmquad3xpiperxmarginrescmd;
wire [1:0] ifpscpmquad0xpiperxmarginreqlanenum;
wire [1:0] ifpscpmquad0xpiperxmarginreslanenum;
wire [1:0] ifpscpmquad1xpiperxmarginreqlanenum;
wire [1:0] ifpscpmquad1xpiperxmarginreslanenum;
wire [1:0] ifpscpmquad2xpiperxmarginreqlanenum;
wire [1:0] ifpscpmquad2xpiperxmarginreslanenum;
wire [1:0] ifpscpmquad3xpiperxmarginreqlanenum;
wire [1:0] ifpscpmquad3xpiperxmarginreslanenum;
wire [7:0] ifpscpmquad0xpiperxmarginreqpayload;
wire [7:0] ifpscpmquad0xpiperxmarginrespayload;
wire [7:0] ifpscpmquad1xpiperxmarginreqpayload;
wire [7:0] ifpscpmquad1xpiperxmarginrespayload;
wire [7:0] ifpscpmquad2xpiperxmarginreqpayload;
wire [7:0] ifpscpmquad2xpiperxmarginrespayload;
wire [7:0] ifpscpmquad3xpiperxmarginreqpayload;
wire [7:0] ifpscpmquad3xpiperxmarginrespayload;

wire q0porresetn;
wire q0sysrst1n;
wire q0sysrst2n;
wire q0sysrst3n;
wire q1porresetn;
wire q1sysrst1n;
wire q1sysrst2n;
wire q1sysrst3n;
wire q2porresetn;
wire q2sysrst1n;
wire q2sysrst2n;
wire q2sysrst3n;
wire q3porresetn;
wire q3sysrst1n;
wire q3sysrst2n;
wire q3sysrst3n;

wire [552:0] unusedtiehigh;

wire cpmoscclkdiv2;

wire [14:0] ifbufgtq0clkbufgt;
wire [14:0] ifbufgtq1clkbufgt;
wire [14:0] ifbufgtq2clkbufgt;
wire [14:0] ifbufgtq3clkbufgt;

wire ifdpll0pltstden;
wire ifdpll0pltstdwe;
wire ifdpll0pltstrst;
wire ifdpll0pltstdclk;
wire[15:0] ifdpll0pltstdi;
wire [6:0] ifdpll0pltstdaddr;

wire ifdpll1pltstden;
wire ifdpll1pltstdwe;
wire ifdpll1pltstrst;
wire ifdpll1pltstdclk;
wire[15:0] ifdpll1pltstdi;
wire [6:0] ifdpll1pltstdaddr;

wire ifpscpmcfgaxibuser;
wire ifpscpmcfgaxirlast;
wire ifpscpmcfgaxiwlast;
wire ifpscpmcfgaxiarlock;
wire ifpscpmcfgaxiawlock;
wire ifpscpmcfgaxibready;
wire ifpscpmcfgaxibvalid;
wire ifpscpmcfgaxirready;
wire ifpscpmcfgaxirvalid;
wire ifpscpmcfgaxiwready;
wire ifpscpmcfgaxiwvalid;
wire ifpscpmcfgaxiarready;
wire ifpscpmcfgaxiarvalid;
wire ifpscpmcfgaxiawready;
wire ifpscpmcfgaxiawvalid;
wire [15:0] ifpscpmcfgaxibid;
wire [15:0] ifpscpmcfgaxirid;
wire [15:0] ifpscpmcfgaxiwid;
wire [15:0] ifpscpmcfgaxiarid;
wire [15:0] ifpscpmcfgaxiawid;
wire [1:0]  ifpscpmcfgaxibresp;
wire [1:0]  ifpscpmcfgaxirresp;
wire [3:0]  ifpscpmcfgaxiarqos;
wire [3:0]  ifpscpmcfgaxiawqos;
wire [3:0]  ifpscpmcfgaxiwstrb;
wire [31:0] ifpscpmcfgaxirdata;
wire [31:0] ifpscpmcfgaxiwdata;
wire [5:0]  ifpscpmcfgaxiruser;
wire [5:0]  ifpscpmcfgaxiwuser;
wire [7:0]  ifpscpmcfgaxiarlen;
wire [7:0]  ifpscpmcfgaxiawlen;
wire [15:0] ifpscpmcfgaxiaruser;
wire [15:0] ifpscpmcfgaxiawuser;
wire [2:0]  ifpscpmcfgaxiarprot;
wire [2:0]  ifpscpmcfgaxiarsize;
wire [2:0]  ifpscpmcfgaxiawprot;
wire [2:0]  ifpscpmcfgaxiawsize;
wire [63:0] ifpscpmcfgaxiaraddr;
wire [63:0] ifpscpmcfgaxiawaddr;
wire [1:0]  ifpscpmcfgaxiarburst;
wire [1:0]  ifpscpmcfgaxiawburst;
wire [3:0]  ifpscpmcfgaxiarcache;
wire [3:0]  ifpscpmcfgaxiawcache;
wire [3:0]  ifpscpmcfgaxiarregion;
wire [3:0]  ifpscpmcfgaxiawregion;

wire ifpscpmchannel0xpipetxswing;
wire ifpscpmchannel0xpipetxdeemph;
wire ifpscpmchannel0xpiperxpolarity;
wire ifpscpmchannel0xpipetxelecidle;
wire ifpscpmchannel0xpipetxdatavalid;
wire ifpscpmchannel0xpipetxcompliance;
wire ifpscpmchannel0xpipetxstartblock;
wire ifpscpmchannel0xpiperxtermination;
wire ifpscpmchannel0xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel0xpipetxdata;
wire [2:0] ifpscpmchannel0xpipetxmargin;
wire [1:0] ifpscpmchannel0xpipepowerdown;
wire [1:0] ifpscpmchannel0xpipetxcharisk;
wire [4:0] ifpscpmchannel0xpipetxprecursor;
wire [1:0] ifpscpmchannel0xpipetxsyncheader;
wire [4:0] ifpscpmchannel0xpipetxpostcursor;
wire [6:0] ifpscpmchannel0xpipetxmaincursor;

wire ifpscpmchannel1xpipetxswing;
wire ifpscpmchannel1xpipetxdeemph;
wire ifpscpmchannel1xpiperxpolarity;
wire ifpscpmchannel1xpipetxelecidle;
wire ifpscpmchannel1xpipetxdatavalid;
wire ifpscpmchannel1xpipetxcompliance;
wire ifpscpmchannel1xpipetxstartblock;
wire ifpscpmchannel1xpiperxtermination;
wire ifpscpmchannel1xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel1xpipetxdata;
wire [2:0] ifpscpmchannel1xpipetxmargin;
wire [1:0] ifpscpmchannel1xpipepowerdown;
wire [1:0] ifpscpmchannel1xpipetxcharisk;
wire [4:0] ifpscpmchannel1xpipetxprecursor;
wire [1:0] ifpscpmchannel1xpipetxsyncheader;
wire [4:0] ifpscpmchannel1xpipetxpostcursor;
wire [6:0] ifpscpmchannel1xpipetxmaincursor;

wire ifpscpmchannel2xpipetxswing;
wire ifpscpmchannel2xpipetxdeemph;
wire ifpscpmchannel2xpiperxpolarity;
wire ifpscpmchannel2xpipetxelecidle;
wire ifpscpmchannel2xpipetxdatavalid;
wire ifpscpmchannel2xpipetxcompliance;
wire ifpscpmchannel2xpipetxstartblock;
wire ifpscpmchannel2xpiperxtermination;
wire ifpscpmchannel2xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel2xpipetxdata;
wire [2:0] ifpscpmchannel2xpipetxmargin;
wire [1:0] ifpscpmchannel2xpipepowerdown;
wire [1:0] ifpscpmchannel2xpipetxcharisk;
wire [4:0] ifpscpmchannel2xpipetxprecursor;
wire [1:0] ifpscpmchannel2xpipetxsyncheader;
wire [4:0] ifpscpmchannel2xpipetxpostcursor;
wire [6:0] ifpscpmchannel2xpipetxmaincursor;

wire ifpscpmchannel3xpipetxswing;
wire ifpscpmchannel3xpipetxdeemph;
wire ifpscpmchannel3xpiperxpolarity;
wire ifpscpmchannel3xpipetxelecidle;
wire ifpscpmchannel3xpipetxdatavalid;
wire ifpscpmchannel3xpipetxcompliance;
wire ifpscpmchannel3xpipetxstartblock;
wire ifpscpmchannel3xpiperxtermination;
wire ifpscpmchannel3xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel3xpipetxdata;
wire [2:0] ifpscpmchannel3xpipetxmargin;
wire [1:0] ifpscpmchannel3xpipepowerdown;
wire [1:0] ifpscpmchannel3xpipetxcharisk;
wire [4:0] ifpscpmchannel3xpipetxprecursor;
wire [1:0] ifpscpmchannel3xpipetxsyncheader;
wire [4:0] ifpscpmchannel3xpipetxpostcursor;
wire [6:0] ifpscpmchannel3xpipetxmaincursor;

wire ifpscpmchannel4xpipetxswing;
wire ifpscpmchannel4xpipetxdeemph;
wire ifpscpmchannel4xpiperxpolarity;
wire ifpscpmchannel4xpipetxelecidle;
wire ifpscpmchannel4xpipetxdatavalid;
wire ifpscpmchannel4xpipetxcompliance;
wire ifpscpmchannel4xpipetxstartblock;
wire ifpscpmchannel4xpiperxtermination;
wire ifpscpmchannel4xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel4xpipetxdata;
wire [2:0] ifpscpmchannel4xpipetxmargin;
wire [1:0] ifpscpmchannel4xpipepowerdown;
wire [1:0] ifpscpmchannel4xpipetxcharisk;
wire [4:0] ifpscpmchannel4xpipetxprecursor;
wire [1:0] ifpscpmchannel4xpipetxsyncheader;
wire [4:0] ifpscpmchannel4xpipetxpostcursor;
wire [6:0] ifpscpmchannel4xpipetxmaincursor;

wire ifpscpmchannel5xpipetxswing;
wire ifpscpmchannel5xpipetxdeemph;
wire ifpscpmchannel5xpiperxpolarity;
wire ifpscpmchannel5xpipetxelecidle;
wire ifpscpmchannel5xpipetxdatavalid;
wire ifpscpmchannel5xpipetxcompliance;
wire ifpscpmchannel5xpipetxstartblock;
wire ifpscpmchannel5xpiperxtermination;
wire ifpscpmchannel5xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel5xpipetxdata;
wire [2:0] ifpscpmchannel5xpipetxmargin;
wire [1:0] ifpscpmchannel5xpipepowerdown;
wire [1:0] ifpscpmchannel5xpipetxcharisk;
wire [4:0] ifpscpmchannel5xpipetxprecursor;
wire [1:0] ifpscpmchannel5xpipetxsyncheader;
wire [4:0] ifpscpmchannel5xpipetxpostcursor;
wire [6:0] ifpscpmchannel5xpipetxmaincursor;

wire ifpscpmchannel6xpipetxswing;
wire ifpscpmchannel6xpipetxdeemph;
wire ifpscpmchannel6xpiperxpolarity;
wire ifpscpmchannel6xpipetxelecidle;
wire ifpscpmchannel6xpipetxdatavalid;
wire ifpscpmchannel6xpipetxcompliance;
wire ifpscpmchannel6xpipetxstartblock;
wire ifpscpmchannel6xpiperxtermination;
wire ifpscpmchannel6xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel6xpipetxdata;
wire [2:0] ifpscpmchannel6xpipetxmargin;
wire [1:0] ifpscpmchannel6xpipepowerdown;
wire [1:0] ifpscpmchannel6xpipetxcharisk;
wire [4:0] ifpscpmchannel6xpipetxprecursor;
wire [1:0] ifpscpmchannel6xpipetxsyncheader;
wire [4:0] ifpscpmchannel6xpipetxpostcursor;
wire [6:0] ifpscpmchannel6xpipetxmaincursor;

wire ifpscpmchannel7xpipetxswing;
wire ifpscpmchannel7xpipetxdeemph;
wire ifpscpmchannel7xpiperxpolarity;
wire ifpscpmchannel7xpipetxelecidle;
wire ifpscpmchannel7xpipetxdatavalid;
wire ifpscpmchannel7xpipetxcompliance;
wire ifpscpmchannel7xpipetxstartblock;
wire ifpscpmchannel7xpiperxtermination;
wire ifpscpmchannel7xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel7xpipetxdata;
wire [2:0] ifpscpmchannel7xpipetxmargin;
wire [1:0] ifpscpmchannel7xpipepowerdown;
wire [1:0] ifpscpmchannel7xpipetxcharisk;
wire [4:0] ifpscpmchannel7xpipetxprecursor;
wire [1:0] ifpscpmchannel7xpipetxsyncheader;
wire [4:0] ifpscpmchannel7xpipetxpostcursor;
wire [6:0] ifpscpmchannel7xpipetxmaincursor;

wire ifpscpmchannel8xpipetxswing;
wire ifpscpmchannel8xpipetxdeemph;
wire ifpscpmchannel8xpiperxpolarity;
wire ifpscpmchannel8xpipetxelecidle;
wire ifpscpmchannel8xpipetxdatavalid;
wire ifpscpmchannel8xpipetxcompliance;
wire ifpscpmchannel8xpipetxstartblock;
wire ifpscpmchannel8xpiperxtermination;
wire ifpscpmchannel8xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel8xpipetxdata;
wire [2:0] ifpscpmchannel8xpipetxmargin;
wire [1:0] ifpscpmchannel8xpipepowerdown;
wire [1:0] ifpscpmchannel8xpipetxcharisk;
wire [4:0] ifpscpmchannel8xpipetxprecursor;
wire [1:0] ifpscpmchannel8xpipetxsyncheader;
wire [4:0] ifpscpmchannel8xpipetxpostcursor;
wire [6:0] ifpscpmchannel8xpipetxmaincursor;

wire ifpscpmchannel9xpipetxswing;
wire ifpscpmchannel9xpipetxdeemph;
wire ifpscpmchannel9xpiperxpolarity;
wire ifpscpmchannel9xpipetxelecidle;
wire ifpscpmchannel9xpipetxdatavalid;
wire ifpscpmchannel9xpipetxcompliance;
wire ifpscpmchannel9xpipetxstartblock;
wire ifpscpmchannel9xpiperxtermination;
wire ifpscpmchannel9xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel9xpipetxdata;
wire [2:0] ifpscpmchannel9xpipetxmargin;
wire [1:0] ifpscpmchannel9xpipepowerdown;
wire [1:0] ifpscpmchannel9xpipetxcharisk;
wire [4:0] ifpscpmchannel9xpipetxprecursor;
wire [1:0] ifpscpmchannel9xpipetxsyncheader;
wire [4:0] ifpscpmchannel9xpipetxpostcursor;
wire [6:0] ifpscpmchannel9xpipetxmaincursor;

wire ifpscpmchannel10xpipetxswing;
wire ifpscpmchannel10xpipetxdeemph;
wire ifpscpmchannel10xpiperxpolarity;
wire ifpscpmchannel10xpipetxelecidle;
wire ifpscpmchannel10xpipetxdatavalid;
wire ifpscpmchannel10xpipetxcompliance;
wire ifpscpmchannel10xpipetxstartblock;
wire ifpscpmchannel10xpiperxtermination;
wire ifpscpmchannel10xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel10xpipetxdata;
wire [2:0] ifpscpmchannel10xpipetxmargin;
wire [1:0] ifpscpmchannel10xpipepowerdown;
wire [1:0] ifpscpmchannel10xpipetxcharisk;
wire [4:0] ifpscpmchannel10xpipetxprecursor;
wire [1:0] ifpscpmchannel10xpipetxsyncheader;
wire [4:0] ifpscpmchannel10xpipetxpostcursor;
wire [6:0] ifpscpmchannel10xpipetxmaincursor;

wire ifpscpmchannel11xpipetxswing;
wire ifpscpmchannel11xpipetxdeemph;
wire ifpscpmchannel11xpiperxpolarity;
wire ifpscpmchannel11xpipetxelecidle;
wire ifpscpmchannel11xpipetxdatavalid;
wire ifpscpmchannel11xpipetxcompliance;
wire ifpscpmchannel11xpipetxstartblock;
wire ifpscpmchannel11xpiperxtermination;
wire ifpscpmchannel11xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel11xpipetxdata;
wire [2:0] ifpscpmchannel11xpipetxmargin;
wire [1:0] ifpscpmchannel11xpipepowerdown;
wire [1:0] ifpscpmchannel11xpipetxcharisk;
wire [4:0] ifpscpmchannel11xpipetxprecursor;
wire [1:0] ifpscpmchannel11xpipetxsyncheader;
wire [4:0] ifpscpmchannel11xpipetxpostcursor;
wire [6:0] ifpscpmchannel11xpipetxmaincursor;

wire ifpscpmchannel12xpipetxswing;
wire ifpscpmchannel12xpipetxdeemph;
wire ifpscpmchannel12xpiperxpolarity;
wire ifpscpmchannel12xpipetxelecidle;
wire ifpscpmchannel12xpipetxdatavalid;
wire ifpscpmchannel12xpipetxcompliance;
wire ifpscpmchannel12xpipetxstartblock;
wire ifpscpmchannel12xpiperxtermination;
wire ifpscpmchannel12xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel12xpipetxdata;
wire [2:0] ifpscpmchannel12xpipetxmargin;
wire [1:0] ifpscpmchannel12xpipepowerdown;
wire [1:0] ifpscpmchannel12xpipetxcharisk;
wire [4:0] ifpscpmchannel12xpipetxprecursor;
wire [1:0] ifpscpmchannel12xpipetxsyncheader;
wire [4:0] ifpscpmchannel12xpipetxpostcursor;
wire [6:0] ifpscpmchannel12xpipetxmaincursor;

wire ifpscpmchannel13xpipetxswing;
wire ifpscpmchannel13xpipetxdeemph;
wire ifpscpmchannel13xpiperxpolarity;
wire ifpscpmchannel13xpipetxelecidle;
wire ifpscpmchannel13xpipetxdatavalid;
wire ifpscpmchannel13xpipetxcompliance;
wire ifpscpmchannel13xpipetxstartblock;
wire ifpscpmchannel13xpiperxtermination;
wire ifpscpmchannel13xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel13xpipetxdata;
wire [2:0] ifpscpmchannel13xpipetxmargin;
wire [1:0] ifpscpmchannel13xpipepowerdown;
wire [1:0] ifpscpmchannel13xpipetxcharisk;
wire [4:0] ifpscpmchannel13xpipetxprecursor;
wire [1:0] ifpscpmchannel13xpipetxsyncheader;
wire [4:0] ifpscpmchannel13xpipetxpostcursor;
wire [6:0] ifpscpmchannel13xpipetxmaincursor;

wire ifpscpmchannel14xpipetxswing;
wire ifpscpmchannel14xpipetxdeemph;
wire ifpscpmchannel14xpiperxpolarity;
wire ifpscpmchannel14xpipetxelecidle;
wire ifpscpmchannel14xpipetxdatavalid;
wire ifpscpmchannel14xpipetxcompliance;
wire ifpscpmchannel14xpipetxstartblock;
wire ifpscpmchannel14xpiperxtermination;
wire ifpscpmchannel14xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel14xpipetxdata;
wire [2:0] ifpscpmchannel14xpipetxmargin;
wire [1:0] ifpscpmchannel14xpipepowerdown;
wire [1:0] ifpscpmchannel14xpipetxcharisk;
wire [4:0] ifpscpmchannel14xpipetxprecursor;
wire [1:0] ifpscpmchannel14xpipetxsyncheader;
wire [4:0] ifpscpmchannel14xpipetxpostcursor;
wire [6:0] ifpscpmchannel14xpipetxmaincursor;

wire ifpscpmchannel15xpipetxswing;
wire ifpscpmchannel15xpipetxdeemph;
wire ifpscpmchannel15xpiperxpolarity;
wire ifpscpmchannel15xpipetxelecidle;
wire ifpscpmchannel15xpipetxdatavalid;
wire ifpscpmchannel15xpipetxcompliance;
wire ifpscpmchannel15xpipetxstartblock;
wire ifpscpmchannel15xpiperxtermination;
wire ifpscpmchannel15xpipetxdetectrxloopback;

wire[31:0] ifpscpmchannel15xpipetxdata;
wire [2:0] ifpscpmchannel15xpipetxmargin;
wire [1:0] ifpscpmchannel15xpipepowerdown;
wire [1:0] ifpscpmchannel15xpipetxcharisk;
wire [4:0] ifpscpmchannel15xpipetxprecursor;
wire [1:0] ifpscpmchannel15xpipetxsyncheader;
wire [4:0] ifpscpmchannel15xpipetxpostcursor;
wire [6:0] ifpscpmchannel15xpipetxmaincursor;


wire ifpscpmlink0xpipegtpipeclk;
wire ifpscpmlink1xpipegtpipeclk;
wire ifpscpmlink0xpipepcieperstn;
wire ifpscpmlink1xpipepcieperstn;
wire ifpscpmhsdplinkxpipegtrxusrclk;
wire ifpscpmintquadxpipephyreadyfrbot;
wire ifpscpmhsdpchannel0xpiperxpcsreset;
wire ifpscpmhsdpchannel1xpiperxpcsreset;
wire ifpscpmhsdpchannel2xpiperxpcsreset;
wire ifpscpmlink0xpipepcielinkreachtarget;
wire ifpscpmlink1xpipepcielinkreachtarget;
wire ifpscpmhsdpchannel0xpiperxgearboxslip;
wire ifpscpmhsdpchannel1xpiperxgearboxslip;
wire ifpscpmhsdpchannel2xpiperxgearboxslip;
wire ifpscpmlink0xpipephyesmadaptationsave;
wire ifpscpmlink1xpipephyesmadaptationsave;

wire [2:0] ifpscpmlink0xpipepiperate;
wire [2:0] ifpscpmlink1xpipepiperate;
wire [5:0] ifpscpmlink0xpipepcieltssmstate;
wire [5:0] ifpscpmlink1xpipepcieltssmstate;
wire [1:0] ifpscpmhsdpchannel0xpipetxheader;
wire [1:0] ifpscpmhsdpchannel1xpipetxheader;
wire [1:0] ifpscpmhsdpchannel2xpipetxheader;
wire [6:0] ifpscpmhsdpchannel0xpipetxsequence;
wire [6:0] ifpscpmhsdpchannel1xpipetxsequence;
wire [6:0] ifpscpmhsdpchannel2xpipetxsequence;

wire ifpscpmpcieaxibready;
wire ifpscpmpcieaxibvalid;
wire ifpscpmpcieaxirready;
wire ifpscpmpcieaxirvalid;
wire ifpscpmpcieaxiwready;
wire ifpscpmpcieaxiwvalid;
wire ifpscpmpcieaxiarready;
wire ifpscpmpcieaxiarvalid;
wire ifpscpmpcieaxiawready;
wire ifpscpmpcieaxiawvalid;
wire [15:0] ifpscpmpcieaxibid;
wire [15:0] ifpscpmpcieaxirid;
wire [15:0] ifpscpmpcieaxiwid;
wire [15:0] ifpscpmpcieaxiarid;
wire [15:0] ifpscpmpcieaxiawid;
wire [0:0]  ifpscpmpcieaxirlast;
wire [0:0]  ifpscpmpcieaxiwlast;
wire [1:0]  ifpscpmpcieaxibresp;
wire [1:0]  ifpscpmpcieaxirresp;
wire [15:0] ifpscpmpcieaxibuser;
wire [15:0] ifpscpmpcieaxiwstrb;
wire [16:0] ifpscpmpcieaxiruser;
wire [16:0] ifpscpmpcieaxiwuser;
wire [3:0]  ifpscpmpcieaxiarqos;
wire [3:0]  ifpscpmpcieaxiawqos;
wire [7:0]  ifpscpmpcieaxiarlen;
wire [7:0]  ifpscpmpcieaxiawlen;
wire[127:0] ifpscpmpcieaxirdata;
wire[127:0] ifpscpmpcieaxiwdata;
wire [0:0]  ifpscpmpcieaxiarlock;
wire [0:0]  ifpscpmpcieaxiawlock;
wire [17:0] ifpscpmpcieaxiaruser;
wire [17:0] ifpscpmpcieaxiawuser;
wire [2:0]  ifpscpmpcieaxiarprot;
wire [2:0]  ifpscpmpcieaxiarsize;
wire [2:0]  ifpscpmpcieaxiawprot;
wire [2:0]  ifpscpmpcieaxiawsize;
wire [63:0] ifpscpmpcieaxiaraddr;
wire [63:0] ifpscpmpcieaxiawaddr;
wire [1:0]  ifpscpmpcieaxiarburst;
wire [1:0]  ifpscpmpcieaxiawburst;
wire [3:0]  ifpscpmpcieaxiarcache;
wire [3:0]  ifpscpmpcieaxiawcache;
wire [3:0]  ifpscpmpcieaxiarregion;
wire [3:0]  ifpscpmpcieaxiawregion;

wire ifpscpmpcsrpcrapben;
wire ifpscpmpcsrpcrpwrdn;
wire ifpscpmpcsrpcrmemclr;
wire ifpscpmpcsrpcrgatereg;
wire ifpscpmpcsrpcrscanclr;
wire ifpscpmpcsrpcrfabricen;
wire ifpscpmpcsrpcrstartcal;
wire ifpscpmpcsrpcrtristate;
wire ifpscpmpcsrpcrdisnpiclk;
wire ifpscpmpcsrpcrholdstate;
wire ifpscpmpcsrpcrinitstate;
wire ifpscpmpcsrpcrpcomplete;
wire ifpscpmpcsrpcrstartbisr;
wire [3:0] ifpscpmpcsrpcrodisable;

wire lpdcpm5porn;
wire lpdcpmtopswclk;
wire lpdcpminrefclk;
wire lpd_cpm5_por_n_int;
wire lpdcpmswitchtimeoutcnt;

wire plcpm5irq0;
wire plcpm5irq1;
wire plcpm5refclk;
wire plcpm5axi0clk;
wire plcpm5axi1clk;
wire plcpm5chi0clk;
wire plcpm5chi1clk;
wire q0npiclkepxpipe;
wire q1npiclkepxpipe;
wire q2npiclkepxpipe;
wire q3npiclkepxpipe;

wire [31:0] plcpm5gpi0;
wire [31:0] plcpm5gpi1;

//q0 to q1 connections
wire [3:0] rxpisouthin_to_rxpsouthout_q1;
wire [3:0] txpisouthin_to_txpsouthout_q1;
wire [5:0] pipenorthoutq0_to_pipenorthinq1;
wire [3:0] rxpinorthout_q0_to_rxpinorthin_q1;
wire [3:0] txpinorthout_q0_to_txpinorthin_q1;
wire [5:0] pipesouthin_q0_to_pipesouthout_q1;
wire [1:0] resetdone_northout_q0_to_resetdone_northin_q1;
wire [1:0] resetdone_southin_q0_to_resetdone_southout_q1;

//q1 to q2 connections
wire [5:0] pipenorthoutq1_to_pipenorthinq2;
wire [3:0] rxpisouthin_q1_to_rxpsouthout_q2;
wire [3:0] txpisouthin_q1_to_txpsouthout_q2;
wire [3:0] rxpinorthout_q1_to_rxpinorthin_q2;
wire [3:0] txpinorthout_q1_to_txpinorthin_q2;
wire [5:0] pipesouthin_q1_to_pipesouthout_q2;
wire [1:0] resetdone_northout_q1_to_resetdone_northin_q2;
wire [1:0] resetdone_southin_q1_to_resetdone_southout_q2;

//q2 to q3 connections
wire [5:0] pipenorthoutq2_to_pipenorthinq3;
wire [3:0] rxpisouthin_q2_to_rxpsouthout_q3;
wire [3:0] txpisouthin_q2_to_txpsouthout_q3;
wire [3:0] rxpinorthout_q2_to_rxpinorthin_q3;
wire [3:0] txpinorthout_q2_to_txpinorthin_q3;
wire [5:0] pipesouthin_q2_to_pipesouthout_q3;
wire [1:0] resetdone_northout_q2_to_resetdone_northin_q3;
wire [1:0] resetdone_southin_q2_to_resetdone_southout_q3;

wire m_axi0_pl_buser_int;
wire m_axi0_pl_rlast_int;
wire m_axi0_pl_bvalid_int;
wire m_axi0_pl_rvalid_int;
wire m_axi0_pl_wready_int;
wire m_axi0_pl_arready_int;
wire m_axi0_pl_awready_int;
wire [15:0] m_axi0_pl_bid_int;
wire [15:0] m_axi0_pl_rid_int;
wire [1:0]  m_axi0_pl_bresp_int;
wire [1:0]  m_axi0_pl_rresp_int;
wire [63:0] m_axi0_pl_ruser_odd;
wire [63:0] m_axi0_pl_wuser_odd;
wire[127:0] m_axi0_pl_ruser_int;
wire[511:0] m_axi0_pl_rdata_int;

wire m_axi1_pl_buser_int;
wire m_axi1_pl_rlast_int;
wire m_axi1_pl_bvalid_int;
wire m_axi1_pl_rvalid_int;
wire m_axi1_pl_wready_int;
wire m_axi1_pl_arready_int;
wire m_axi1_pl_awready_int;
wire [15:0] m_axi1_pl_bid_int;
wire [15:0] m_axi1_pl_rid_int;
wire [1:0]  m_axi1_pl_bresp_int;
wire [1:0]  m_axi1_pl_rresp_int;
wire [63:0] m_axi1_pl_ruser_odd;
wire [63:0] m_axi1_pl_wuser_odd;
wire[127:0] m_axi1_pl_ruser_int;
wire[511:0] m_axi1_pl_rdata_int;

wire ifplcpm5botgtypfti64dmonitorclk;
wire ifplcpm5topgtypfti64dmonitorclk;
wire ifplcpm5botgtypfti64dmonfiforeset;
wire ifplcpm5topgtypfti64dmonfiforeset;
wire [63:0] ifplcpm5botgtypfti64dmonitorout;
wire [63:0] ifplcpm5topgtypfti64dmonitorout;

wire q0_ch0_rxpkdet;
wire q0_ch1_rxpkdet;
wire q0_ch2_rxpkdet;
wire q0_ch3_rxpkdet;
wire q0_ch0_rxoutclk;
wire q0_ch0_txoutclk;
wire q0_ch1_rxoutclk;
wire q0_ch1_txoutclk;
wire q0_ch2_rxoutclk;
wire q0_ch2_txoutclk;
wire q0_ch3_rxoutclk;
wire q0_ch3_txoutclk;
wire q0_ch0_rxbyterealign;
wire q0_ch1_rxbyterealign;
wire q0_ch2_rxbyterealign;
wire q0_ch3_rxbyterealign;
wire q0_ch0_dmonitoroutclk;
wire q0_ch1_dmonitoroutclk;
wire q0_ch2_dmonitoroutclk;
wire q0_ch3_dmonitoroutclk;

wire q1_ch0_rxpkdet;
wire q1_ch1_rxpkdet;
wire q1_ch2_rxpkdet;
wire q1_ch3_rxpkdet;
wire q1_ch0_rxoutclk;
wire q1_ch0_txoutclk;
wire q1_ch1_rxoutclk;
wire q1_ch1_txoutclk;
wire q1_ch2_rxoutclk;
wire q1_ch2_txoutclk;
wire q1_ch3_rxoutclk;
wire q1_ch3_txoutclk;
wire q1_ch0_rxbyterealign;
wire q1_ch1_rxbyterealign;
wire q1_ch2_rxbyterealign;
wire q1_ch3_rxbyterealign;
wire q1_ch0_dmonitoroutclk;
wire q1_ch1_dmonitoroutclk;
wire q1_ch2_dmonitoroutclk;
wire q1_ch3_dmonitoroutclk;

wire q2_ch0_rxpkdet;
wire q2_ch1_rxpkdet;
wire q2_ch2_rxpkdet;
wire q2_ch3_rxpkdet;
wire q2_ch0_rxoutclk;
wire q2_ch0_txoutclk;
wire q2_ch1_rxoutclk;
wire q2_ch1_txoutclk;
wire q2_ch2_rxoutclk;
wire q2_ch2_txoutclk;
wire q2_ch3_rxoutclk;
wire q2_ch3_txoutclk;
wire q2_ch0_rxbyterealign;
wire q2_ch1_rxbyterealign;
wire q2_ch2_rxbyterealign;
wire q2_ch3_rxbyterealign;
wire q2_ch0_dmonitoroutclk;
wire q2_ch1_dmonitoroutclk;
wire q2_ch2_dmonitoroutclk;
wire q2_ch3_dmonitoroutclk;

wire q3_ch0_rxpkdet;
wire q3_ch1_rxpkdet;
wire q3_ch2_rxpkdet;
wire q3_ch3_rxpkdet;
wire q3_ch0_rxoutclk;
wire q3_ch0_txoutclk;
wire q3_ch1_rxoutclk;
wire q3_ch1_txoutclk;
wire q3_ch2_rxoutclk;
wire q3_ch2_txoutclk;
wire q3_ch3_rxoutclk;
wire q3_ch3_txoutclk;
wire q3_ch0_rxbyterealign;
wire q3_ch1_rxbyterealign;
wire q3_ch2_rxbyterealign;
wire q3_ch3_rxbyterealign;
wire q3_ch0_dmonitoroutclk;
wire q3_ch1_dmonitoroutclk;
wire q3_ch2_dmonitoroutclk;
wire q3_ch3_dmonitoroutclk;

wire [7:0] pcie0_s_axis_cc_tready_int;
wire [7:0] pcie0_s_axis_rq_tready_int;
wire [7:0] pcie1_s_axis_cc_tready_int;
wire [7:0] pcie1_s_axis_rq_tready_int;

wire pcie0_user_clk_fb;
wire pcie1_user_clk_fb;

assign pcie0_s_axis_cc_tready = pcie0_s_axis_cc_tready_int[0];
assign pcie0_s_axis_rq_tready = pcie0_s_axis_rq_tready_int[0];
assign pcie1_s_axis_cc_tready = pcie1_s_axis_cc_tready_int[0];
assign pcie1_s_axis_rq_tready = pcie1_s_axis_rq_tready_int[0];
