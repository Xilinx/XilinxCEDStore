`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Y3LVj5yZZiI22L0qPUFDZF3JNAKSietZHuiC9m5WO9ijq60ilfX80y4PLp1+Vfs2TnKWKoc0gs9W
mXUXlgM3z6ysQtsuQ8GG4dqazDNvStgsPgeb7guHylNEN2w6cX/HdYWl/LH001osG1Adkx83Vujp
f0WBi3eJfirdOn/n+pJEcZytNdmyX3N/rJxu693vOUsS229FQ0dUYp92L7mxORrKChrCkwxed3xo
26LVRSyjhhTUxAnCNAhEi923kfwNcFyxqaUQ7+FhAth9mio56qSJP8+fIKnD4KqO9voiCMjHUhcR
aEkpPfX/gCiezyEKHVaJsJE+AjCFFwt1g4w55g==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
RL4cGExkroBpvGDDclPJ8InQ4famJpSctpjOR2O/G+LQ5xsrntkiAvWwmQB+E8lbP3AAwcs89dMD
fU7MqC8N9YZH7TVN16LoWwo7TZT9PzBlcLZidetLHiV3ANQUj+tcD8zomF7jfMFuz+snxWTCLsiA
NrTP3drwh+Y+Bm++BA9YbR6xYByKgDuSD5MIng+QEstoe9LeJfzIE4EkKyOhHd4gGfgWCzOefqft
pEbNhHdtRU3wqfglohhbqDnq37roGl0eAvbPGONKM8CVCb1BzahsxlDkeGiVA+Kc+68HZx/+Pllq
NQQLJ+6jyYBXhmsa4NiF5sSQoRAeYGdds83LBGQw1tR5Mm81AfmlinPtfnoX1aGmd63SUwdqJTey
tcI04mLyKMcUNNlqxdoQFP+rc3+OYmiFJh4AtF8CxlaRAicFKbBA1niLO3G/ZnYqAOS/mslK6cz2
a8p03FFK0qncHB99daIAnXSENBQKJIjso4wd7Dl+jMwtwz42/o4PARyR26TufTZoyhdsRSqC3HAS
kRru8e1ACiWiVONZVfS/qduFnToK7TcYS6pDCYMcudWyagyJdsTQ0WBPOCiHPzyde8TUbvHuUKjB
ZRVjA8mon94eEOGblMabqOU2Z9Nteo/w68zAPeb/zyABqs54ITYU4bClRMmJ2j/gyqdQe+kSojBK
APz6bIsrvJzTi3ZgZkQfuBFNIUMDndscPDwy89j7b9844byDKaI6VgxZ9jd2Q4hzN07P/878cu3q
OffFAvOrQRpyjmwUPjO2ZmyIKdjkdGD9f5sD1YswDqWhEBy7Q7njWCIxMIsyhTk/Wu30hfu9iEBP
DwvANeq3aQxH6nBSXiDMa2zuIJ539DOSQOEkoRTb4oW+tw4zg7ojGpH6UvTGRpsqKiD4ZnjHz5xX
+OTvBCaAXmTKh4dhb2710QIZm4d5MdvgIIsVqkM43cZM9UVfMbTAiMqtwiYtld/g4Mxac62TC2rn
7ala4BNPZRptuU58k4NskYssnjXeZRBJo6JCxUXRFUtnSoUJ4G6K/NHX3xhBozny+2vau4B5qHz9
HsBqRieDiwqJgP6Gq2kU7cQi2i2b0w0+getxiA/30tUt62TCPSkQYi4UVJBkXEH1G2n+9UKCavEM
u4daeaxuHeknd0Pcarx+dascvSPeIFgzEuOOb9eUrpj20NnYSqio3HAOLbvo04KMO1IkTF5tUBJR
gdd+fMPlQShuIU2zFAgn9Y1rl5VV4T7b9/Qmp+qcIoU9IpNUe0kJTqAF5vIjkdTVz7OtIj/YLTYs
C9ISAlmxwncn3tXQRU5Yagkb/IeGPgi/gND5EXm8big7bJIXKSFkZElaAwzgxqxIfhAQXImEVIIY
m8OalnxlgCqkTlT0tweQC0WGP8De8C9hguN5mTA3yuEg3q3d5Dt6FnqWCo8CSQR/ANGpPkRRhT9Y
NgxXaPKPhfejRnv9mL55OryvzhKAGD7K1O0YdN8dBlzof0ty2NphL8ZQuwEDdu9Lehb+ETLLJpnb
0JR3Rcohbs0QjbHqnmZZzpzkgdeYMXiw0mIgU1TqCiLZsZYyjcYBHjX6NnzE8kyyXKnEndFqFntp
avTzt4ZXJTf16zK+hYtmbMSEf8y0baRFIQW9EfehyHoSTThmNybw8l54hhMrkW8OkDQpoXEbOsOq
63SC50qFC/mwwDTPzCiIP964DENxZAxE4Oy+FH//jkCQPII+bDgm9TByTO+nbZ4S8t0X1uGcHnOz
Zf8RIdU/Hz3M2Ae1kqyQUsekIsGpn3EEmKMz9uyQGF6sJNYH/7YOtuo8YHY2u2zsTAviNbodcfL1
tffLloq9xlbSzbacRDuH6ahSURuplmFVJwFD/5Og7hI+6zlNIEEA38Y+Y6vY791h7glg3Q4fcNaG
nvN924xOtHrbcgLqN5Xwms4dyGQTGBj51jWSz1GFvDu0GyUq5kEI4MRiSsNeZwZXvCDlIJ4WN4Xj
iupnjlcxqprVkPB3ix/qMkGzZKdHH5Js3ds4GY3pYIuQxUxKOe2B5iI748sgdY1v1KS+KSPvuXun
uDXnh23bBltSaTrohRej+E570ozyvArBptcdO+3iHdZbRGOM7JxOi2pvW2EYPJHSoCVLvIEEFtB6
3Tmrzui772El+MC/cZiDymZMBlMqI0oBRYQKemCsYRnohHeVzflLbpYgw5rIA5mBBi52CYqVRb6X
ATVn5AskMrQ9JubU4LcuSWGv49Gs+9y+446iMQMHlE18NrKP4FNEr/MXaUBIqW4KqbmOK20Sttpx
idj4dQPEKtbMGNuUNP+e43fpL+TnDIt+mhBK0riN3lG8vB2KvBMRjbP+6C+WOxWAem0X8z1JXc6o
Z6ixbEG2Z3/9CxMtXkTxFif3PLusR5bf0EmWEjyeRXPfFQ5E2h9Bzxg6XKEh9ZaIIIe6Q7mN6Fht
DPlrGPwzjIBC5S5YP1bGDk+GMaRlVyPwAzwOyjdJ2ejee0Yh+COYKNtvfAUSqlI1ycGr2SqfsgP5
RmFox8PolsvDPRcmpNUYcI/veBdg4kFohFsTq3vyo4c3Y237dFYlW6/n4cabI+cposMd8Cy9rWBo
hxVwENa+lhtD7PK7up0B7O6WTuTlgAdnqNAsEv1nI5BSrRRrDJ+XpjnFaxXJX4guMka89vghWj6F
roRIbuWPJ+YpSFVG9jmawJ+0kdcmZEcrDs7oqWM8wUtD9NU6CIJ2ZnpURryh88kKkGi+KZT+U4Bq
ownAIHaSBlxVmDLEOKH/0KqXjXUazNKYegUD+gadao/CLy86kPZmNZqwsj1HCypxvtJKiPElGz4W
oLko6guodLKG1YY1UoZnreiuErxkocJ8fdZF5yUVeo+OsaFkyK/w6CMc5kkrHweg1qbEUwkqmVhQ
5SDwT7YyfU2guzfW84QJsUWxNymbrheyfFLJNidQ2i7wse/MzWMvKwuZnjvFIyRInOcEH43kKZGf
0tqplgsV7UUamQOavohBuKfqC57LcvbPalVoEdO8GoJGWcRj+mt/rLPNKvL3GenpG/iFQ4HWt8/8
T2ch1guzV8wZrFj4lrqUumhKKTzWq8qBQxbHzFHJZynNWtQCH3++RYPUposX1ktza73CjepspMb8
AkQ7txTHrk3em2OpuTUU1jYtgQJSHJmUWMPGiEc01edEccmIZSjw4z5FQzbdfDkeAgN3nlAySKFP
3aFyDGkUca/x43kELWFqrewACfGXQ0qx2RbHXEfFwNwaoXjDFphQWbju+IIRUWznGUQXBU68pKPe
zmW5EI6k/5EIlG3YhQ/U3MAVCJvAXU/sjN+PfPAyg93pm24m+1f0aKL0JgoWXmpdz5n0u4Kb6s75
tUyts6/klVLIpJJ6bdiWvLnVo78cf73onKO4ez7qXdQN7QK33mtt9sfJgo9xCrQVSKW2ZOL7gp41
e/TqIHb+Eo0YnymvFVAWGRplyFLjzcH7gL92tFUDqvXp8fTwrtqgmtWzdqfN5bn6PNfQwGzez1GC
4tSP8eXOOwUGmW/LYhyuTRSTJWDyW0Y8bVVvNPlUhCcyfo0KNpa2u9zSoeYFlE2PYKcTaaV8RwPa
7HzdTCqt6SEvod57wEHGkeVyMAiKVFMnOQNeh5KJyrUHGTpBEG6NPsHqwHKvCcCdQtEAAegh1JRi
OrPtkmcPqTP5rU9XCDpAbR3tE1yvJP2RZhxQRok52xbox66tIIooBZjfS62mvXWNfV6PUZeL2RRT
MtflxdDSm2HKq0OM17dLMsCFMU58jM6GEpmSXQMhwmv0H8eb0nLncO8wDTt+O9SM9Xff+mKLxov9
su5Ajfih+Gbyq3fiPMmOwqODIxT0ZpaTNHViv53ODiNJ03Y7J0nrxUaqki8BWvJfdK8/SQl138bn
1lB/DT7j+QEVOTuSRR0GTn7sdyPYaM7NKCwvdK13vM+2bezA1ZC3TjzTbfKWMZeQf5qvbPQkut5J
+ge3zDQGCzQtuXLcKpPwGfnkNiRBYbX9aZFCU92vivFukP6TAkAwpquYFqt7MRg0P/ETfYt6tIH+
lYYSbo5GwdN5r9Ie+WdcKGuwoBOiQCrDSxMPykaypxxBFOggh5KiBHhMMaFhsoQOSAQJG84s96pn
RLuKD4yhONrbAFF8HWM3nd0cyNRsKwS75F+2EQd0JVlPtgSiYY3m38GzbATxTyPnhnc1dl7a/c9Z
hK6U2FV67ay6RS/Ft6P0VQW5VAP7CNNBLcxpPHVZK9O8iCFSbF29sGLmxrP2boTFbzlhZ/QYrQi7
cMoQnaBvSol43B3f+r8DpSNIUUvVf68s7gtZXffFD7Po95qiSWjy5ur9ej0YXck/6ILG2gdkaAQn
N4sxmGfOzzX/gQNQgnSvSqSpA5Ah9hXCMv6kc8KsFy2iDu+KNGAHhgnRsQEHcPxuzRlqVRXW3Hk1
EU9PFvJ7hnC/H+KCl+Bs5njdjurPPmc6rdiv4S/hVthD0tAigfiKTQhK3BWxUWFVQImyE27XQknv
5RkkT572qdD8QXo8awwTl4oM87Aai+0sZDUQ93Sa1OwivcwdOnecEYFDjWpHWgiqbeWAHWeUsIhz
YPw39825GNAJZr78c9JSabCFRHzIdKx/KBPYzR8cdYdkppp2ISP+jLUwxihlXqBrOf5abrfXmFuY
aRVH9UL+17zPrDe62YfKrBI8XUIlnTxFiLBBx8C8mQmHmPNPdhmor3gFY5CktgFfJIqXrdawHpEp
SNcukA6r24+eX6qHDvseB75iO9OgnZss65fu4E+YUpQZdHphZQq7FAb2IgJgEKAPL4EtgimLCZZa
Z8elItteX5I16BEIG4r8SUGV/lnA43WcZmn/197hu+6iZX0wxWTrft1ExWTMnX7DePQOfTJuJExI
EQqkpioh4kvwzFkO83QIkTehAW7Wd16GxaGgpP98elWJW7oPbPwjT91zHXOhznczK7MMKAMvtV9e
OYNTZI6I2T/FZ+kkAdBL9V7hykBxGeVqvH7B8tITuV5N1ySe5lMd5RNQ3DFOFL1YeVES/s/M3+YF
aPOnb9RGHh7p/zojA6MpheMVmST5aywx3wsn+xjuV3YCivRdf2HDmCz1byRBcUT9AmaClfAJPbRG
ybp31Q88jZyQtoidmcauJhXNYFuBwh/SbLaGfjx/het5rU+GjZztzihpuDJpXytj/moKZPEcFVRb
7voa4WwTTBbqd0QKB1/FIEHTE4mysixMS2lyic6EV19vHqH6R4TRefO8w0ZUdft/7NN1EE+w4e5h
MP1aOqVcgfJov3FeUhn53DXXMe0sTCH9dMlvXDjllocYKrYShf6EpiTNoMqelmn+gZqnma41LtFS
7sfjP4P/E4VqLtfRGqp2i+J8KhHIK6VGTPflS/F2hqi5YkrTUe7KUrnYNDcaIC8Scr6IWYJykt/B
ceSDVqfe4KdK/Zbg+kg/vmilJvKDOppq5bb6D0eq0eyC90jPdka99GN5GAy4FQqaQYh9BM1KOaDZ
fKQg29lIg54aYIP1Q27kUFIuYZ19/C9S2Z0wrvgZ0iZMoYgyqvLjySS0DWe9BH1S/UU0kOXvup2A
JLWzgbzToYjCpeO4QyPOrnZ9aVSMuR1jk/levzTk27EsDOUgAs0To2tPrAz0P+pOnorfqcrY3kI8
oQ65sg9DwtJubsWCO6WEZWPwCJ+oRVqDkfB4DbGJaZ0u32nwirDXeiVPQWO33OKkCd0CapAYqttP
EmPFTtA3HP6E2pUK9wwtcZlODEBlQgXIHexyq7Ud2qT3KTqu3IrW6ODw5YVKg1sWqKrWK06pAATA
pziAe0C6g7RqAAjfohLR8F2FRObmOl3rHQ41wQFs90Quov8sXneXsCGR6hGNZwYbRmoS4JlbAi4p
axHwZ0Z1kfZN20Yyv2eSsTXDrPSV1dBSbt85jp2xIorP4kfQjSGqBxIm5/XLIGicWqK4AgCXbfrV
D2JiX+wXyGbX43t/hP4vwhMeyi/ToCB7Y37rlIGz14fWytEvzC2wmOeK+joOs9FzyqYess02FGM/
H8yFP3KSVeWJeN9/5LQ5HuUqYeNdAeVnZiTWQXWIId7ABkwfXXTCyPCbb/Q+31CJJIiIHVrlDpek
LxRNmzJ76J+S4ovk0n1qI7FUw9VhWq6fGRtvEkjZqCs4BlbbdHoK2q+L2tb38OJ4Pe+43vmXPnqm
7anSNpG3kJB/KeZeL6REAgDKi60ptXJrprRq5NzRhgdbV54M4nxSw77nAKz29MnH19rweDe7SaAX
a/azHolfHRnDuzrliZmiKZcGN/6h6hXxMFHWBG8wzS9J2ONVRJa3GLiHJg/Hr5g5PUQuHIt3Ce4i
qBMMopCm2UbNPyIw1CakSGSIeI7e8GCDB0yjh6Kt59/R2KmWlNXicQ0vCY3CDusDLZ9giU9tQby0
bMOx4xIeVl20vNP52x1q8YS8UsUjiQKhGHtRjSopK0dB39gxFKulTN3NndpqTU2QaGDBPjSgXRj0
hGchq3oycdjDFXzy8Ui7XtDd93pRRZqn1UyYVniXVVtv+aNtOEQRpq1tdFPq+HR0RkRkkSwYgp/p
othgTqw+4tX+fCUaC5Sx+dFiT4bVWIg1nG/THA7jxRDtlVDEwc+/APCh6pYxnEX4+GV2FQljGX9d
9onafdPYKSn4lCLhbeVidgdXCCy+wDlJsl/BPwNIPUFBvjMu9toYu1NFX/NCZBJKdAlf0tgMQNS3
xEfJPJbpQH1URctNOO84DghEoid82ulujQvRK35sA7vI+k0XY7W9/XiNVg02q4fWpnitp9fK6Itv
Nl8P/67JtBlwyi5X2B3hAaaVNtqKXrdao6IptjnabTinlRsTgud+qenUV+HnJhkKZTrt6GcjE2ig
pW3yijJBEPnkMgJGLumb7IxuKbHWal1lEzNQQ7cMPP6SNUWlnNX35OFfEQPR7MLXohkp6a4hZBzM
sfIuoe9qX3UXd/ASf1+ONGyDn/eTB2gN7Nvd2wsC3Gszg/IspdGTqVXmka1XzYwPqiElGjT06zCZ
cUNMPENJvYVp0usZh2zbcZIWNqlZHEhJo/7CybE3KbzM0sX2gnHQXz2wCLkkoqexYusBhmOp5fD7
Ns6su2sJF8hSEIH/fc8tHwy0RyOg0J1WdJw/zY7a0czbohvxtw5LqGev8wCx6QUraVsoJlPvCsIO
PN9jM+aSvyHWW3RoUcEeT0nOn5BMeaykP0Zwel2k8oyoF/3ufxJNF0ZCiikv0OQF2QUAlz3cB09B
9Q2yPCXYMEkEHmEccw+3vxxgoZduRVbQtzJH2klWhITv8gaMOlWt6ikcxJ3C9Xc02R8OazkpVdzR
cqpKSnMjIJl3y6v82yGQVnmKta3/QC/EGwMJaS41Shcv/ao60cLVaj9vib3FczLlTBcrbWs3V+oy
Hw7ynC39EUW5OlyNHZor1mbhcpML4debgVbUTEnuwGQbGenqF2zjDDu6Tz2QWir60HaKK65KlMrV
d1Kv8/B3j5B+g8c2/iL8REzAzUt7pqBxbDRDel8ji6DUnw4r5Zx7vdzJUYTSpg80BljpMxtRnM7r
y9crW2KHJxIgWyQDOpxHSrK9dFI6GY7tpXVhmC6Nr+rXwwLv5AmNA7Nbs/3tRwBIu1NxkuSFBiX1
0ZFKgrr0gachff6Kxyk8hyspxCnBYCQoVejj14ObC35fBqyYso87BvB1v3FpL1h63YKFr+naDR5O
4a7ZYRDSYaScrGy8sKVzqzuHamFGaTGK8QBjzbqt4KYGNbcuhigrqhJVBhGlLlZ0TSEp0RkSQjpo
/7HlREf0aQplgft3/H9l1aaZ29wJiFgjAcvovfyJiTG8dMvYqLiofPAjG23vjYVgRG98d54jRWgC
8j+ji0PWYsVItXyGUqgJOK18OhX3us6BTzoCc0SztGFsjKTOHk3zKZIeedJn5tl9GkF02b+hZhdx
1IviRd4GDQuL9TIhvfCaypvim1ibIT4UGoTRKyTO3J9zMcOCAN6uRIPoSqqJBhRx7b6PyEphtrHe
4mKxFDBEhSJyxM+hbl4pdHFfqIEle5AgA5E7P/QSTDIaGEOjlLNjB2n4Yh8AHARWkip1NWjeLuKC
ZlEOfSwp4RcvdQY6QP5PNNWnnglCfUn+KaVfyTlsgvFodBfFHhrDt2X6thpqvrLK48UpQrdw2gMa
Kwao7hQCNPbeZ+mqmsRTMYcu9ZWaNoBb5im6zSzpYoPG9UbNm+ptUWCpJpbyd07jnKuW3L/n/TDF
/aQccCxOk1yso5P8qaMI1KFxFmVxS3V/Gx/F67qT1+71yOUOgcJrdzgN8iMoK+IwWWBAHoTqlMzy
6+XqGufe2yGnYHEO59zQKBN51M3VJGZAyJqRK9GbGNaKKHhmCC5kVNTmaZzPoeI8kj/n8r6tYyV4
CIt/pX0M/fstJcKXOFFu1B2VH2josag1EqGyuvFGOeB3TDyy8dMBHWtNrRo6cFVqwrKqhhvPIM1J
Sp96uqtDqGYuMbDdhNOGjYXwIiCPR62eEyypHj2A9/VesbzMMbWTZNdWvHyEDZHEYGzXqV7ru5PO
eVktDbHbasb6zQYkn2usnQVPunubT01DgkT1is40qXYTbpDmW5vlmkhJpVIPIIChXwH68vUPYVcw
VsxCuYJT/KCRS4duHg0GfoGsYqKHYEwqDwzMZhg7lKuJTYhFNvgPyyQELm5OjrSwY15dN+UPt2y2
Z/cq/E/xgFmt6fxxFC2xvoCpcldustKlf0obigH7ulq68DO7IxJkdIIcAD8JgCPYc/sqEGxuEPH7
5MM0Yu/z93h/ZvSpfJ29zHrbKArSKzdGxD4K/yVSLlgus/xT1L6mwNO6b5Yc1G++r5aqy+s5qGl3
5Q2DnYBjkx+NAMGGmjWKCoBcty3eCh1vxvJPvSY3ECi+0h5+w8NsUGEhuGwaZLA8nBXFFHkG5Rpl
kj/JfucCJKKFXH211jesKRmn9idZmBSr7rrdHIyGoV3XPHBXv6uR9whFw6UKK+7R2yJ3CewdqmAf
nv+MeHl7wObwoywbsmNoZzrTpH2tdKWg6xq/v6mGhf4PezQoxicC8iQ8kA2GxEX3n1TgYDUWSnEX
PvvaphhHPzN6agjNrFlXKjSQic9Fcn6q4s8oCTgLEyy0wBodu8B9LKkz4chBErlHUeG4lsxvOtM5
MteC5Fe8dH5gMXS7USBzmh1X12EPG0ezbiJcMaKbr+Kx5hhLWAq2YFzx96j/MI5+4PfnffO2eUS5
APnPinQmm334m73aWbYSJyVPKLZNywSkgWYhNRi9a+ptjN6wbX45AvH/ux5humLhN0cFVmEEWdfP
x+Jmet/PY8F1pQrcO/GEeOByLXy7gq/NIsb5PVf7UD8Ie6/UYBLHfiKw/Llwgs5W9KgkeFrQtkpg
tNjmHgTf08baKiR8flqpBHoZNKpsJDrLGRWiNiUmDjoALCHbvopbFiad6+YLjDzBk7VIP97RAYXB
DGFDQzy/DgQo6Jx4EMXuHo7Byd2uTLSKQmCwa0uXtgN+yW64g0bAuRGOwOshz2XE6l6xDmPeycKm
qB/aGOSu7lSLVxcMrGw7JEjhFdQWfX+vnGcPlK+/ehCD9v9SlKtKsWdbQpPQis2vKS2H/w49V7xy
lq3l4e7PrSskuQQGizTxwllTJR5jEQNsfe0LTGZ4BtXEcfumCb8p1RW2/twkg+uozy9t9IGIu2QM
vAz13iouT4FEPbyIEeCjszjrqlaq1JxpAO/Lf1wxLWMfmSka8EJyNVNOPaywlhB+cKykBSqU4dHW
rGhKUhxg0bBO6RGq683U0rhfnjefx9xQsn/0qDjVXniIXHepV4UZ4pFMTYiSoe1WGfkyjfYNsUgn
JhUxi6dlBKKbpelr+PQo6x+CvKGlXn3yEsSlcKepMl8nq1J9HOraWaB616vcGw9An+TPLTVljzpo
Is19suEpFqO9YZbSs2hq6gqMXaZD/vViCizy+OzTmkLuqWXaOm6P0aOigoAJm95ua0qaESzVxCti
mULTK/EkS+pfD4qxo3MrV6ZTkXVNDu60/T8q1Dt2Cq/ns6JcfPbGcyBVDhw9gTW3a0Z0ppfRAxdn
K4K3uMZdWdVAhCimG5uSICFznY+DBEBkSUAn7Pov0BcaQa3Xbw6rAG8URDqycwh/nAYtkVGuTYHH
X5lZD4QSxH4FptqvKwNZjhcHoJMrlRP+bQ+eEEp0ttRF31mGBR8xgFfyaTOjzsNlX4vE3oDEvz6e
a+R1yiISixT+hWwrCDHpz1em0yW6LxPyOErkyc/dcMDlw6wau9UQUeriECcuKWRBpC1r2eH/UMgv
x8aXWGuTAABPH62Xi9W5/4WrRDo2M0CyKYf41zSnVzT8sKahRVi95YzQh4ZRjJ9631dOMzcRG064
hox+UxKhbDb32MfT6ShsoxtmF0T3Xiq9bRlaaEefSaA7B1EJKivsTGXH+p2Myfuxi7a9cl22EXcK
N+8OVpuuXo9T884speXOPCsj+1DOF2ojHXFPh1lCkhjElLgZDQleX6TABSZhAOHMl45aB/xwg6v3
95nKwpT1j6G01oD4oBWwO/GVfzd2VPDffWllzIDaYIvz+UGFDexCgylfdnAcUtBECLRJdcW04dwQ
+uJ0lUNfKzpeyqKu6hZ5JZLyBIx5U9NJB4EqvVWHkRKa82YDlTjuHAHkSG6jLVeqmeGv92NelvLP
fFipA+iU/DhJO05qNlrvJHyDVdJpHHPtaomWarKSyBuPmuFPYagT2GhdOMyeTdBEk4qUT9Ul1hkw
DqJ71WVhIGfRRv3oaMkNBSUk2sKil1WNPUfE+lBeX9OADZWgQV3qz9h/ZIE//MnkPqz3DLBTccRT
psaB0pIZ989Yb6ikZZ2BDAnmGKv3ZbyBvAoXzVCyl9d/8bZd7cP4GWr3hi0PnRf/PBjEmyzZ1RJq
QomDUNtuBquK5Kda0URVyhy069UbPdU8oWMKJkVU4PlRTaDXI+FrNtoVQ9KUcw34VQDUvERdthel
R4zsc77J/WB2nfhhxwNJIeyN+sqlwlCTwxYuGpnmVWevMY1MDOZt4Bby5DeU7uNW2dF8LEKUwYZS
iucmAnxOiJbiSziAFGcAYWR74WuZsZz9oCqn3bAB/Pk7kufAfkl0/5Z9v7BMCoeesEt/UnpX0iRJ
tsXE87CTIrwl1ff0vbb1fg2vCS5MMkvuUhXvjZuTnVGnvoKigixrl3X+FjHPJryNuB2M5pHZ3k1V
leqRLCJM909vneOxt4tR0f6qxEZj+A7juMd3pyq/n6PI4VzyUtJjuDeXtIAX7pkvmwMdTt/dp24B
LhUXL3NQ/Jjjf33CnLR84ly3VNqr/oLEprbQpcd76S2XGGVVQNFIjhNCJ5WU2XsZaOyqUo5QG3z2
0gKs1A3priBNFsvwbFKYK1qntHayydWjwq9ZUi8t7CdxOInNO0AF+QIGuo60slsi2ZCUdwUfU8EM
I+0aLCP0b5eRGUnepRCwyBUbZxYrCKcPJixT2vuNwqURUwrJggNFGBPcOn3hG146MO4KQKxkkaf+
NJWezaAKJyxXPdt/ettNpVKoBjonjYqmBJpOsCfANTJZJUydF3skQREpxFC4WSYMEbY5bE2YRI6O
5eJJa5DcLSjJ5ZS7EXtPuQTMzDfnHJBovki+lUW2EfdTUui7we3lEZxVDT2jSK3MusHtpiThzKCM
RgSQaGEQ7OAJDQeeEQ/bDF6fPDSLHrtfYbO49F9iieAquKr62IKIXrLf0ydoQz5WwilX86ZMMmmR
K08qTlJw5vgz+acYfLd4XAe80okZjYH+lCwL5Iuah8/77XcF2DnFIArJoXbevRa5mvpUFm9g9CGo
uHN0ucHpjfuKLw5ph6gRMvYrufXe73NoqLYBKZKZ+aHSkkinijN1RKbaqpg5WpYxqXnX1x1/TkSc
+XSKms9Mw25akGTdZTqgI8ubKGpah49ga88MBbhf/qPqyYtn/TtSwO8X/nU3mj6OqFA1s6P3pX9F
R9RvHqSCW/xdCtnJZVZnY5dxah7aS3BvUT7j2wqC6pas9MS3ZlvRAwb4JAd9k21h22wsdgsA22xp
nF1jKgkU5Q33yb1XfIK7YVUYgF5/tN9p5vHzwxTL6gdiiiWzQrKkEqu/cYbDLkDSxppfoePnwiwc
+1KcLfkhgV2CXs02II95KRLBJNoopfpdwB38Ett2dvCJQaBXiLaperx9YBN2vGIig0Rzgf+cP5vc
L+01ZQypkBpjb3oXG+6yQK40bmPPyPZ0n2C8bj0iFGSkIwOHmPvNb+3ZcUvvWde84ZZUAydBw1XU
N+NIftNILDgi8xObkkYjBTo9il4Zy713rESP/wkHWWmlLrmX6YJwVjV6AQ9HWhqGlCDLZDroKxOS
nw1CJ2Igqfw89Fs1EvCuhT2tcH8jnxNa3xZZ9M9KBWcbfSLvfwWCpvTj3wMg943JLKISyNrMsTAh
tQCDi2So7mNGJ3Vre+vqoCgBM7BMrItO0BWjmv/AnSYXMo6EajLUwsgupUAc7xbREVuWPAKGizHQ
7b8pUYr869tPFxFD/A9lTGF6+6SoHLO8cOcJwJWzHSueUFesDOEitlYGTsfvKhWZnDLL57CuyQCc
PJahUKED7ap50pZ3dmtuAtuYJ0wF/hFNPiVUsMryuxR1jPcGsdnymyNOafaBcDp6czDKoHnDSTqj
cN28nHujFyf2HF/z6vqOCcGxRGTeKdO/MaEwc9TSacmr/tfwzkalvHGJQm/DoUDtQX+/PZxsHpp3
+UjsWlnlclHqXtGytc2GI5CUtofl24xfC5rF7hkVPsx6rMopevj94CRSnTSAoLS01gw6r3eqoalY
Pvaxa6CB/sw1qJG/j+ZSJ2JWPRc1tzriwnFxfpsXwXmsmy0gqyBnPu8q9w6HOyBr82afEXVnw7ZK
3DaVA4jTGMAI0XFb1KwirU4IG51sYQST9q+P/4w+EjdxN68HZkhm1rOms31jdsvQtfSQVUITq48u
RDPsh3O86S6IFwkP85J6/cMDvpeCqpj0choVco1mt8mHAHiFKcDJjtxE+jck5CY987LxGSPjr86v
DzZKPunfhEjc3fDY9TX3NocDV0euaEeU55gbnxc/8CuUurPCRbZDNGVPbjlA4pb/RvL4TMA5FoWH
8e7jHXj4zmDVTDhSnCLVraCoh/Q9jUEtXuJhMPTmxTWYGoyhOk5ViLHoWL2u1FX49700E46OQVRq
01u7K1rhdi8uwGFQ42XXUYXcg7JkWxtQ8WDWw2Aqy6YwOlIjqmfxDxvvgvwcis30i9CyzAYJ+gvj
2W6xBo9aesW8pyf0rBqdonyVJ5Nsv1HFDTvMLczBjnnunSFlXv+bGxKKVtPQJAhAJl50JUPLJked
JVnCT61J4MqzrsSWxpwSZg+VCz8qSEYUqHcsDLKFMiIg9u19FN2UBAXub6MM3zmPTTNBSugCdMaG
N0RvU1TF69kpilL5RoYRZ+4biRXehzJHm0UzbQJXsSYgAFLiwKJwRpHeJcH7h0nKr1Oi29+Ch/NZ
gZ4hLDhajONuG2+9cghitXVqWZBUZx6EGyJ0jeJvjc9mjaPDGnRPRt7vzFBTbNDe/WlwP82faGEP
ukz/DfEVNsSz8UrsI0bGzhOTfvTOGn8uAeI96H77GwBp69Ss8+7svBlSMM9HGr7n21WyvbQGZW0I
DfcJTU6CGk4PXpSFk87rM3IIHwPUrLZ0cpNDpyqJ6mAbJuy38sw6cQDO24/yXYFAPhCW+kJEgZMz
84Zk+YGHHMfib7z0VGo0n1LFZRhRJKiAtiMKDbfEpk/oqkZu4S3KWqgOVtkhA/ggtNRy6ULo8USh
FRPIH65rQoXqIsvqBQdAVyp1GfC4HyMW0lb3z/Ib6XiI2xwCP+FxVQNpAS1qqHvoFnCdUJe5uASp
tN0jX4PE3rMhILQmYllmlRaJA9u9HMPGYGhU/VGHtY5VHlmEp0hV3SkCJJz4/Hgie6cA7pK9bsCb
fU1iANJ+BOw7hMLd0bvWDlqqJ+sX2hRq8vX+ToYr82b9CEWkqeSkuqbzAvBCPb/C+AFVE3WxhRmH
nvYRKXut9ehOeUkAbXkI2kFjn3GzLmPJ+ubsmLvn6b10fiXoQmOoKcg9OlBsKeKzZ2BflH7yo18l
kk9kBMp/GlR6vT4lvWbEkiq7gKWQ0MsnVFHMfaN73O7aOcw3cPKbM0hEMvzR9vKIaFknMthAeICv
SZAfBOTIzu0SSUDDbT2ShsxD+cg+4ckxsd+yHqhXOPJLGofb9kn4vWFNLNbp3uipYjhuqJkRMuaq
ATHeD7gj3OG1Q2HCaFxRqsiTkwtrqVmJ0o5G5scdI6SW1PLn07o6mshbzrcn6OuH0KvkIA4yGboQ
RvCnwEqc/5T1yHx+0QfzdPXQQO7ftUHGcPjWVh4vMFwzw9KHvd9qw8kn1hllhTBUqhjPQSy3nGCV
iLN9217UBt/TfOrAXePOpT/ap5TMsCs13Q5jI3eOAF1qpEbU5J+YC+BSHRa/Xnu70cnw4MyC3Ur6
MO0a7eWUzoVncssCupsTqGZV/vIaCO0JSoFnzUIG9ASh4+K46db5IV76aRkSGZz5ix0Cmt2hMtgb
Udf6P7WbNLySKHqRaVocgzC7lAK6P+UOA4/mOr5De87P26dTqY5bSXF1LFq/2FHUQgfFzlFeTjuV
17O6LDmKwwXoDqS/fYjmcB5zv/6XqI/DefmEgTREQQGmpd+M3BBuW1A40pxn1g2bcBOcJlcYhHFf
FDpNlSKe3otm/NDt+9tuqe3a/xpDeG0ykqXO4KfgBZSMsIAPEVaBUk/76swH9HnIJFo3R1PpSMuL
I3EVaNP/D4yWbKOyKgeep8VBD5AraEtuPF+yn/5uKwexjpRmHF33QS97VGLh/jW4cLP8afC42LkQ
LQPwQbfePNyRUVcwD0UWfDO4VXz7GtZRzhxnSIlJfocAnCC9Ahuo0ISz9LAwAMhyWzxi3mz9u9TQ
Qnv4/3KLP/wWZxNcXs8pKLr5JgVSLlAIr0aoM+uoNeOImIvJtjVjgYhILXs1KJNbl7TzrypDhpgi
gOkmxdxUo87JaXWsdRuTLOkvLCuPsduTLfgg4SzHJNUTvEsbsI3Yb75V148DxQjVTEIjUPKdRBMZ
OdovFLrC0JZvGVOHhgcK3NKhAEaz2JpnWKYjmxeDn/A02Zv0lzGlmuaVK6pN8hBmP970PZRJxWvt
LezsoR3ySMKXjqViPoX39bHKz2eAvtVLn/ZIN/frqVEq/ez7lWOqjr5KcD0PdC5n2TEK2Mer3Unb
b67azWa605bXcsT/xsup+lfx9ixKZbhYS8ZR2BZULi7GqaKOU7u8Lk1+jQhghbmP9XP9I5wVDypJ
cNbDtD+mwVXk/DKWZtsOcqfL4S4EHzu1LwMVUuDjyGLrFCtxw84Jme3Fk/zJ9kIx7xZ4Yf4FRxnk
Q5j7ZcIheTHwkrE6pBT/ECfwYzL/kaLOvJRDDMvf3SyxfH7wGPhawiaJaofEKGsno8uvlfunovX5
FutLoHm+MmkbSgijk3y+JgoxcHzShIjoZlYCCs8yyJueE3qlyD6v+0Kb729KkRwhzGllW35aEr6X
3JKXON0LKm1jHPLYzfzLb/OCoDDvO/qkMzy1v3/b6Kk83YAwE9dCpRN9jcW5oomwT7vCa+2BSSnJ
EXClrVxHoG8hIPMHI1LaLvVjpNsiaMB4y2HfMdeTUe6cLfUb0TUH3hX/pLdSNBiP1yJxAvByqqAr
NvT+Cb/67ccBOVMoBL9k0ICGZcbgzj222fHBR1UYS0GE+yZGvFN+OZha3Q/QSG+Ho5SZahDbN8B0
mIMbhc5Ij4BJjjxxRhjSanVHtscuzZkbMb1y8nvpBD+30xKunxrF4yD/hPDHN2mZiKu0wgAxerfA
AaQv35HnH5kwXqO57qplakkBWBGt32bgtJo0yjRR8iMWBp7baSziphX7OcIlWB/X4ksd2w867uUj
0pnoWkvWpPWAjm6gFGBLDzbQTajBwkpY0ddmaIbA1w//Uyg+N9SRYbQ4wJ8DLIwJBqTOBrAUg6+z
nyXf/nOPMpHSrRPMNS0qwTIOnhJmeIL8qOw6elC6YExTfOwMxW2ddqsr8HY4govStSrp3fIjLK2L
Hwdve/+YpA7Jz2fahHVMXYQSHs1ku0Y/7uAg+r035zjc8p+x0nRejKIvRjOhVM58WHot5Lk8ns3L
iPctvTFOaxQQmiqEa+FMQaTdSVZ8tipLuh5uMo22dZs7+u8kLFLHZqVPsUIneE7w2xkZck5W7cOP
6wsx8kWcTjwscX3Kpx4D6t7IuBuWwOgbnQ5UbtrNI8LOn/PbL5NpXhj9GCusl5oWCt+X/lCEbzYH
1O5rgTAyZDvsIhK8CwjZ1nPNB3dKDPPASlfot74Hrp6j7829kgc6ATT0eLNL43DpCn5ouyoqXlmC
+HiNXy8799/IWoAeuhjmZZdbZx9EUt9cja0xrTCxygOHYKwgbbt88avpQoWfcyFvQuOneKPGr6pZ
+JHsJPQpk5CfI2wwnw6QIbV6845IlEdYdHdtpothb10t4dAl/YzMY/4bViTky/8CTfq2JMggdNI6
fxynBwzjeMbniCFfolZhtBUEiFN8AwQNcSCBPE3hrtXMBVUdQzqR1Jc3UYBlFBrd1709Yr3pNKaA
+Hhdk0NQPqsezfUq43do/zDl3wb+I2PFB//KEDpAz8TosH1m2QRFk3QSpY3LgNkGW8NTpv35RR/b
KcH9UrQsaHW2XhVsoHYIlMhmyovzJQ9T1TFHRZaPVxCVMYD405pOC/kHRcTE9xVu7WukhQd/wNQO
tH9OZNuIrNedohNs3w2V7deYXcVzNSTCq7wUlHiDb1y6UHC+vuJuqp9kTkL5PXumzf78dplHoyea
KbKldoKMYAz8PrY2nzUiDx+hsvcNzz+LMKpOwO3+Sso6wVYe4DXFwUcMxORNQLd0vlMrUZ7ARxzL
J7aastBvF0B97JuZp095HS8mqx7iRV/M9EqE9PGIy5SMqgnTqcYUK6Uaglt7TXGzmOAst9Y3EBVt
QnMH7Ay05nDTYPU2RWv4CGLtOsdHjMNSsbom0u+odTyeEWpSh5VO9syH/0AH3Eb8GEE9nt8lOOhG
qQQ7x5HNIni1CLDtN/aPw7AtEtzMII5U4JYw5APyxrA8pjx4+fIIa1Gda5eZQrT7jN0CvNwX+etr
g1CVEYvwHOCMainobQ6S6o5gWJp7B74eYvWStcWZSsVcYtLPMN9ggHnV2rg6mBb/MDeJMOaYS4ak
KpVHUdq2420vylKsplixMTZ1zGRc1GsKZVcTyQy1gbSef1AQLR/IcLhQBl+HALSeGUlz0H5r6jvI
Qcz+Q6T96U9lNqU9eUfwyOYIEP6nzDVFLaxk7U8kxNYRGWVMIqzolKvFyc3R6+8tUor49nB9ydI9
HhKZgYJ7dq2HXFfLej4Q5SLfM/rYMsSonS1J9wHQEzQzMBVj1i/MQuApfJJy7Gh0Ap+pwChv9xsR
dzXFKh1aoCvxrwGBBn41t/xcwacwpyRft5ieMwjBvR0v3uTykcNWoLNuks/XKKqfWG4faulPusJh
iVsMo121Y7jdSYnearXCPZiX7WTwUTQxjds2DobMgX+dYktrgO8sstzm8tKaLr5XnuVIe97XQj40
kwLhvvncFlcHapNV4/PgGUJJDFRuYQcj2P35iGKY+SAATmQcbRIgJSvHm2WbPDHtJvp8ESaRfXg8
6IZI0sx5kkQ6CyIlymNF1FrEeSQwqIMll+Ecm23PVrBuPQpMAEUBCyQzwaykc08mbICDP85CXdTH
KSGstk33B7iBkFhvoIVcCMqQluiSdCfRm8Y7F5hE+m5sd9oDxJOoEbhEJ9XzLC0mNsoncXHnS1S5
zsxMeByM77tirDJ6zhFDHGNIyZrQsyO9hRmMMBZSiWNC9tx2YrvR7Oq1H1pzPeKqSJDs39kcsGM+
U+yfvfBbXfnmC80c59W4EqKdBjPBhX2kHzkdTvVwQ8b0f1mYoyGeLyyjejIprIK6/YVgFK6bre9J
DqYTnAjnjSH/l8zX6y+aqjk+b1DQc7vrvzBVZO15FMwN1OkGrHi6g35gVunjWecmytAquOPlVfFn
7EenFoKSieRFl15tJABbmaktE0rV3XTxiZjy9GsJ2yEvqSDNb1k5tS2T6ulnk1WGKQhP7nVrUPJT
rbVsdmCDUz6QIkW09zcX1cnqI3HCNBzoI8EArlFmMR773SqRbBAlDwU5M9rppJz4zk8nAs1AkGXV
gHT8YzR8FrqMDnCpq6Yr2FvBSndALVFQyJJiU9DnAiZeGKcvbE8s/gLuy8XwGq1cwZGqoHKO3eSY
zXK7f7CY3vKpCvwH0Hmp87nAHbFr72DVJl7/Srb5LDjRWYEEi1wpWL8YhDPlgyd6wmyXaB6BhL5U
Cbpet1kxfYLNgRO9paKah/CVQ8tA1+eBUDlvA5C0MFQ2XaNfJVznCO/5G5sXsEzf8Vbl7qleD8Ur
CxN7cEVednlZpNn8o+T/R9Xsjs0CMZdqOZZcuf6ZFzenC90symw/NhPDCsdfsqHTipMTHY09mBsj
6K0n34dCJ7xsLd0wOooL2jFsuJSWi9uaByEBZH7Xeuqm/KE4gFMILhXhjr6+6UNzFejk4Jpx8k2V
WXpmr9uxOAzjEgGZbUpM5NXGkJaCsY32+YTNwt5gCYU41r+YPFYIb7ajZf7LUXd1Tk0Ce4FKlhmN
w7N/NrsHezM+NJ1udZWZ3N0XxsIsCDwWSrbrWIBWjcEuARtAz0lcn4/fDma+/1iBZC6lZNMjYg0o
l0lMGNIVH2QIawhoW6fnibveet1Y4w4l8Cx1BouqxFdPbgYktPjQJTXsEOhqFQpfogN/4wUQMpQk
Hb4vIsJiSdVokhQvw8WIIsLuG2UbcpwT6cx0ZnXcbR0GunwBJsdOa3y8HtNY1bD5UdAuWhfJS1AQ
InHjAi0tVzBYO+GHung3O64D7v0yn7VVOJmTDVYOIKvIT0Yc63xsiBuEBmxoBCcxxVdLMKJ+IFoy
rO52wAx3w9eUhZdw5QFdI51hSnA5lKIGvvA+Z0MqSLtrFMyIIBFQdLJI9S7Ym8v3kCuUOJOs3Kvr
BmjWq08CYAkiOTtSICM1L7nxT5LuYIOcyq50QyxjBTliDZzUTf2b11O5Md/JQikeuGQKxnVQKjUE
hqP7XQzz8ldWU1b5n94SyxMLJvlizExbkKGIJmrxs4m2O0by9wpyMhRbwEbQKqYNV5WdapDp09jR
t7mB5w7OCztBy9KSKmSJEHXCcH4aRb2HDzqA17JimJVWIbC3VRSd+tiEN7UxIywXRiQQyZW6rEod
ZWZPE/1hac7KQO1/LI7q480m+1IQ3VoFH/FD4sq7c+5aqYr0lR1tsUig2Kt0z8EGg8/IZkADiCL+
F5jlxKTZLcrtKi7LL2ExH8VCPLS6Nt75OdngG2IkQibdMdxcNyA7E9caad63bEgoEcHE52hPFq5T
veRJ25+rGibCTex9A+fbIvN8mawcpTFvX1OqHQXF8sCPqnBYZ/UADoYUS1pNjM24Edmmg9Xo6svS
AOkUlsnRtOJTyeD/e5CHnKZO7XzRlEHNArsSmEGIJ+u3LJugNdpXvYA13fm6CcT1xo5/ZIZ+xzvr
xEzBYD7VLa2Tv7D4zXUqTcCrqqm304cHQ5Q3ULG7ES6arHhqubweSb22kCyg6HCZng7R1n9ma18G
l8DYrBn0domu++51Rq9TUAh4vX2ZrU666jCdUj27LK+3u+YJBYmSeFWWnnU8nE0AViXRWDfnpV1F
tsAtDRVyh4gWjxJK1QoPJWBaSskbNbDETv04tgBl3PaeczNL1hH8cm+uu1iMfkrJl9AarF7PDlD6
0flEeey/fjG9xTZsUQ/LrE1/vA0wwmLGNHl4udbVfIYmfDw8ouwbO8XqnpNCxacXx2GmGCrWZ+QQ
JHjyNOppVGyOrwijdrlbMwR6g6tl5VAXrW4EVQmxGxcnZCp5Lg3Qz+tmOEdEhQm4gDf7fqsBxLVq
NxBpWgtTkxAXbS8lSQkEkMHeqkWrPPvk3k5QhAAITKp1iSVjQQQhDk5qtAUyzQaBG4HuYH/kWpL8
G/WxKtga7TYXTHsiLWErs+Hf5FTF8b4yPyCzAHAIylurtFefCCoME0dqAEDctW1oY9FCp7OdMk/f
OpPZsI4mG1IIpk4YjsBtpS/gIUCDt81w22AvBMtWMjpIR6b0FyHMWxEtRTIgOcJEUlCI7lvLsxPp
nS5YQos3Neuh2ek0VWyfkjiIR0vIxV7TcuUfhIHqir+pX2kkkneQzjTqkyChImuO389hkFcjyreQ
Icg3BxwVdgxFRtcPSjRQcZz/LQ4s48U5pL0+EwlHpCZK3ZD8GqimvZj/cN2pJQ9SuqQJne3XXdCr
cm9XHLf6E01pbpnhlX6yyyfivwCoXPZpp+Is/xj6q/JkfPFqYBJLaNKXVTZwzvAzYjPqNv9t4rAV
yv6nk/WNV1WoZwMFFdfYI0cJmuNliuldPtaZ4rGTA2B4ukCf9WdrlqJ2011NRG41lcs/o4abO/78
yhEDbk9cFDXWnw05TIOwRi8LRhpWIQakd/sUWTypws2hix41exgpocdKK1UHg3JIpixodLg8xi/n
ZU8J+j/ydyH+Zkj+/XNpDwmJLalCAavXuvB90Rgpr6P4sNP+nI47s4S0IkPI17JVdwqU1RgBgpk4
sIA79MgatHGLDxypkHfgjs0xrlYNenokHDKmCziLPEqFeHSRC3aNHYHSJcW7pKCXh6rmxXo83qvy
i4NkpexRNEDSQmDd+ZaFBfaZ4nJsSu11XC2tl5kUPqkSqbQ2/fu8yDuf632yq/SzBFOaNSR7BAyt
C32Fu5fDVcHm0xJs1LRBoi+/bdRpHYRHfgBKEhiutGpZmgFOBy+mmGJMO9+dSshLkQ1WyVz5vy+j
yxOyzUyh5uiKULoEG1JUEGGvj3BgdOfuPjBYzlkpvAp9o1cXz4sdBqf8AjAenVBO9ii2s/r0nR8l
pvy8TReD5+JMzNYFP91a2uKylKm7IPs8hNiTjI12GDDyGAfWkQU8EKTyJH5ZJEaN1nwHdqgtrzC4
kHgbxAKPMywx4dD7+Cf8zLFnaOMHLYDAHt8r0F0kQR908J3NmCgnkqaH7APaor3OHGIoAuRxZpNy
2+fBprLkSzbb+MhEwv4EbWOuWcYtoVxDexEtqowcwglJ4gk631ZX4FX8T8TD4By5UEDKPjIgaqeE
1M9ItCYzEY0wAAOdDcwsoelGvHiVsqqkYktjEU2CGNsptAJTp7MxVX4w87FVip6BaHjrZtoNcEZ5
VnPo7kyYU07XG42gpl4mGSpGcsR00i4FBA2dJd6QkU2gaT8ezCDg/BczEvAAQF5eunkJSwxWAV87
YBssz0xV4KKk0Aomz74pgwI1LYic59UyoSjQAH/oemayloeU/X+UrQEhzs1bgiCipnBoHZ6WLjWc
m3+yB3DyLbykUsouBGgnpturTVEXpZFeNfi304GEfRQmlj9NwB97iIiuoOdxvqiQfNEK8NlqGZnt
8VHBGm7f+slOO5jG0tZia+XdXKVyrlvWFdiR1bFANPe9M7y1H4HlRen93loXdttSkEP7HRYv6eeB
oXY5yt7buHzHKRFQDZE3Cjg5IYyp1uipvmi0bWBRvVnVzYitEcLsOW9AbhmKkN4ZVegiYkNImvNk
WAmnYwKUkZL3Gz0cIxApxBWi2fQwpgnhJBeLUHcR3m6MbFMZ+HZ10Klc9MHYYgIgEBi3l4pcTGyi
zHSY2qM1n+TmvveTafy0TyFtfYTmJT3iSdWkI0tvYs/de3lW6X/d+Ibu7MnKaFdjYre5jd4UfTVY
XhnNsy5rTBV+nWxQfslGG62dWWQqhMb7Dhuh/e2MvuwNgcsoiJ/tv2zqUMcRc3sQYmb6NptyJP15
RQcESqP4pFeT74VA+ZzAvpipsqWRA1sRFmYbt0/2qN/8swAj9lnAKaH+g2JDRnHIQTlMJrSOhFSt
koFcaqi/FYbE7vMfWJLrJ/dR+k+94GoOELZdkIl/ZQ2XwVfLVDeDst8T6jj0YYn5PJCWgEx9XrtN
nNKByocMpknpKaYdlm6VVkDGMUdPbomUY8R8arR6p1ev7O8ROHDa1vloKdwwQEIowurtJDd6vfSV
0fqIEXiMSGr0Sccxw2mTfb/XILs7C6BGf1LELisGqHpymusEgbm4qEdJecWnY5mH2juVpfxOJPy7
C8Cgl1P9Fpw3OsIPcqlfNmMAV1zU/3Dn0/2tMPtzMOAE6qbYFo8J+0WHoyQqX0E3neh5dqtEM4VH
KEFZLUVzKHUvBXZLGNZ3zGj5Ww6wLoXr7bK7mCc3ve/reYM8R38uh9CQrUj03NC8hhJQAxjJ77UL
3hbReEzDo70joz8qjjG5VRvwwr3LdtNQhT7622ad+21Z4X5+lDPlcpV+S/4wXFBh/l80QllZkCfG
/xXbA+/6Al0eRITaW/ss0I7qI4leQ/8uYOW1CHCZ3dLu8qdLNKKy3l5bu73ZNAxVrmFOysoL/riw
r/+QzZSpWjx9a5B+QMrDrf1JU2kCUI67hFF/BysGWX1fW7Pq4jPVqwdiXMH/QB/Jy+CUqkvDP5q4
rF7dtjfb8zflphxBfI6Iy0cEtl9V5fOBfBdMs9f76EaLOeB9BxneucUFt2JfW+vke3fMi5+aKoBA
icRJb4ScwTKV7KpW+EfiDAaBz8gWRMhnjC3r5rR4P8Q75V4+5IiQP8mLAPYJAbirjW+AHwQtJHo5
HvQ/ILcb45SVWSKH8qkb5JpsrPQ5T64xAxchWMXM3b6hfg1ISnL823WqQf7G2XexsLUSHcEwoZrE
RR+ljLWwPv6qC2hKMWKkb4ZaPKCypz9/mNi/HF++aYy4qGZmS75juF1Aav3A2jljCyVdVujZyA0D
1gQhvFE7LoZ/znvrf10mKo6yvfRTgpVHGHvThp4A/e4egpEFpPpPQEPaJOeoiLH9eZ+xKAAK9CX6
DtoZ5bnRwYYAyV7j6g/ClRGkf8MgNVQSYN0BnuMI4RaJXQOp2rOF0iTSKseA7Giv6DL0TqagOtV0
wxuDo9pOJBbFAJde5Ou3JpETG8n4+VaXR9MSf9076vMj0jTWesyLDcN8wBcv8EgGReJZ0BsFxBvn
zBcE4mMh/AJhfv3JQdiVXkluRIPtvrLdzTob5xq8APHURG92yah2WG1hLLd4tE5vZBm3GBNFwrnW
Vix3jiY2CQRb7WhOJQmUsAobl2vmpPmmPvD3oZXNEme7pxk6Wkzq2GeIv2xuxy36bFjiE2C3sNph
4s1JGpsi+I6qyROSXGWos+HomXtL87oTlGUyNAZQPWy7PX5+IFqUiI9ATLxPdowFa/fUOA2cofsH
BArUTbF7z4WmRrFZBimFuSAWScTy/GIejHNnH0KCiZnx7Wxr00aOv1UcRlszdWAPy0DNQDqERuSH
T5GgZZ6mfT0GMGcI2ehmMxCrVZk9mxVO/62RJNYmuWock/Q9AvGBAhB8wcjh4IL/GiVjqnDcV6I/
V4SKNpK94/8i4ozfU/+Efsihlxgz4cXb+IeDWqGjam/7kp0a+Iu+oAOCpUFn80WiNX/YgkvHP0Tr
XBs8LYr8w4b/HrqHoH4WQkIBF1TfgrACJ+GaLXfinQrvwl6lvaungI0EGHnAiMqZfMSMF3hIQbYs
lfyueWtBWVaKQdvpr9uGyiFtlQZvQFJWzpXdPrhY7aioc9fWDQS92K407JhKaIRMEvw68N3+uOdl
XeqBjjmo0xwipjprdUZ7XMcoU4EAa10NtFv7Gg6c8nhRv9+BmDpJSkRUrVubHFE0PZ2xKR9Nc+WB
cmv+bHMLaulS/GcG6emKr2NkZc3DUFZxSIbs2/Od4evjW74/1cEzKT9aZKQud7RuYsXmiKJEkEXo
xfDWaa/DtMONaBjIRCr/ccfUuvu0Wqb+eJVMD3p8zrPzo1bMgby5bLiX+SOoOdoZL2OPXvHrLms3
egtPm637KxIG7dWzPwjIbSR95wjhCdC+vtcvUsCD0/+A1DAExUfT6BBfhV4eWgZWYCTw7zNR+DT3
YBeew63UX7Bys6Ci860cFfiLEEuI9iBxXBBVG+b0JmoB5gkth39rDap1j3QSjrxu1XcJN59RIPdF
YIIRlXfdMsRrLsoHSL05nfOnO9vXA3tyBopsEVzqpkKZxHx5udX00zPyBIE1P9zpsMvn5X4A8tzU
vayQyRmqfBXA0Ry/xADK3/q2IevYEd8C1MZ9dwT0b9wr9kgDSlMUC4ITavHqrpJ6F4/GiERBqpTo
JAmjlVy2oFQYFUllYCdJ/JC4/KO4BnHh+EdIeAlVZNdw3gdhcOTYdvM+1Hck5st/h2aSb4ZRcwbg
Ty29TskCOzznZwt+De1ox6ghAkkbdq78TDfcu1DR7x/wx9rWHB+P73UtuyaTy2aqW5c0m4MfTMlC
IGZ8pN6L+Pf7iaWuMaahwPMdfRXl7v2f9DXkGfxbjhYz0V/ZDxCJNEOmwL8L/xCUZP9+niMivIQT
4MgKS2yDiXS2i0KzQ8KM1AeRp3Dgk3bPvyzM1w4iLHQCkJmMG84kKg8ylZGgs50X3wMMGVQDlN4D
HTm6ciSeC7mMWAQzYtV8kUaVzFbP573eJkybCWz1/1QZwNlDjjvcbswozuw7x1ba9GkF02cyVIft
poR4BAZ0tIKTT552xvo8clbV5Ehvn1kawbIBzM6p+SGNFbvHq2fNBN+s3iTqrQwUiWZ1uhjQd3gn
roWYfv1a6BPPVS5S8HBbteS3dRPHBSd6WInz6WvtA9kD9r43tz5bsOv31zhCgSxb6q2Yn/gsM7cI
y+bL+jhmkSKax6LpDuLSacI/2lTWNFMIYkdp+pQ7CV9S/38VdNvH8qmtjPqiPFzQvH5MY5qxUIja
i3ertHiA7N//+Yfln6lvu5WxLv7lqEuMx4YDuNCYRMz/RFBfdqVI2jyYOkXHNzXdbcPi0hDBROXF
KLVS+wAD4FvTA22LBEgCABb5ohNnThmjhLO2y3z6Mky93kslr1g+6w11dhchtTxs1uYqhP2Nsntv
g+BnNKprIh7m4KdkbjvJts5JEPKcMNQAtL9jaDWn4Tmbw/X36jaPNpe5NUqIv2XbrfzPtqTB6eXY
K3KVytGbVK3KbpTBwOZjjrz5Gm/FDl1Zp4CahES2dkxTu1q3wo/7x+UwV03P1CP5q4jEg8hErADu
nm7RKYjI+2Adt7bTzo4T3dSIc7tm1c4YoxgALM4DYV9w0b8rzzdq9nrUzfroIIhsx06+59JrqT2W
aEhN5FSV1/n5r18vqC6KK5MenUwmCD61qCm/ahk4a4frWdtH6AhuEn/rnG+HITg6+ofTRLv74uae
6W/kT0+BdDnFPY4lsrGLWzrLcKIhIPD37fmkDNmcHnqfQuTXVArVwGVQyXzRW/1g5jPeSX6dvQHp
7E8GEDjzKLler0sFjqVmhe+I5JhbZGzeVAQzdjJvt4ukKVbM7GYC9e1EQWnwQuoc2wu2U/lmd4ts
rJAmTa7t2nMIuSYsNfNINfwVtXoGkUiMOyIboSL68AuvD33cYm4ZCiWr/9PXRTSo5psL0/yPjtoj
l1IbVnlHYGBvAC9z0/uQAIG1RV/j4aT4PykRES00b7qiW5UCvqP/OyHubvIpk/+UeF4cXqtvFNSg
VSdPJKnytpsB4wbZbrLdR0lyH3+WhSTTl56E++uNAK2utZxwq4vW7CSeM8lkoi6pEtPZsaA2PBZK
X4esT32r77vu/euCMi02pGciz6frC0FWX/OTYBohPfHW6NvPOtW1yhofShUZvWQ8UCgyHyd44TtM
pK8EUJr20Nlur2XZFvmoQtfUNU+QQ19LefYNcOBn2TtxL/0EWFlcnCtaPDgLXozT24unJS4CJEId
N7vTFvK2YaPAxadRhVb0yOkNgxT/XRLGPMQ/qQlhd1bsLrHQcGLGfV/Sm0TuErRzj/a/FzIquOl5
/Rh1Knd7HwDmVHI444Jl9dL/bLWZYX2atXpxYe6TSBLrE+AY/o+RmZcZ3alrMo5MQLYIc7vjVQfC
EM1RQhm0ntnxfcnEoh76xrf8yAkcWOB9tRQ194mPI2u3j9Mht8yhmHy6z7yrM0fNHymKWmlpDYO+
wyXAoPXrhHoyjoW7Z2W7GZbp8dYDA8csXi1xUypYRhsUMK6SFyixusQu/x+ZYnQuVDIFRdie3agB
ngXWLPF/cl0W2AIcosn8pLJVxfTKNcs8j7Ru3h1sVnx8R12WiCIHPYsWVznw/PGsfXYo6zkIHSmF
69mptgojS0FaOGOV7EHewaaYm/4BB+5Bo9V5GrHLJ4Mdim46r5DOOxIXyDe2HZOvnSHTgZiIOsev
NDO9aJc3uNJOgk1tjgbOUPyWBf/lbUjlTGm59VYxto6CqJupIeHlq8/NUGzwISroKZ6G9xcSCCk+
dX0AC/aquqXhrtrE7EKEqwzYE1Ded0N9HZwO53R4jRdoB5he5+SFahi3UpMz3tigBKUrMXHheQQi
/bZ2yEP+uQxD+46lKZO9/UFXbczTuSz2Soz37rPHvN+rkXDSBPVpgXDWZYiD8xdRhq42+d8ViSu0
i1wZT0sVyx/ph1b/uPX8vMlgnoj2dSNG+1Z3BmpJRqilxTWPGh5U2V2LeSh7T5/GBGqiz2eXtrUB
ejxUR0I05K6ArkRUaOjYk28Sep6jydcYYiJVSCa6TdljYJlVZRf7yhEnx8bLZ5F84t3DdWGzEzE5
Fm8fnEo92b/YWxKWWdgzAQzbOtmHG9mJPxOaCqIVRuQsWRqOs4JqD9BWzF2WK+lgvldVkH6fTfOH
en0kKSLMte9OxYUMZ47BQceXU1dEHzx0iOJQvo3NJfnVk7r19wpDn78Lt06WEiZC/L5K8OzLmfBb
r4D+YEw0V9qs0K74aDDE5xQB49U42uJA9qxrDchE96N1tTwmeapYV5rwlnqt14K1grWMITnZxK9O
Mquo1Ce75cUKR84yGc0aQVah666zOmoIBCiDzg1jQPidZjH5AmNr5uFNPlQFxDjIXTY250O3ebx/
wJekg85BXZNG9r26ApCsaoHSIDj3kNjBUagyOZGJavpCeJ7mZPdwrk0yPcOihtwTQ/P2h8dyAOWr
ezcOeRxN0Wu8jxaOkhFTDvqKAlnUy65a33eGXRvetMN5v2yUojY/bp6h9IUHjzvOSQJA+7c2pdFZ
suakoyXua5wNBWCkGOzykxr6kmBhemNFvQpOF1LTAXTjeSjI04Q0wFzP+gnXMdjb+iQCHtMpfREF
xkD17pysnnS/6r4Txpi2+fK1TTXscL0f5wf9p5Puf3RnUIPabmpwHgEkIDR6uabHvLJiMTLkfcSH
mNnabk7bcxXojKbFoTKFGSNx+t0VYibe3gYRpQOs4HrCqV5bXZmlr1bAaZu9jL4ihugpu+Wg4KlU
L4DaLvkXcY+3NRX3p30emv4pLVmslmrn8BLajy23n/3ktYAuFEutbpoEVwxq/zTT0Pug/VxitGWZ
WW6kH4KvHI6KDBOFdInNNu9VPVA4WrOUF2r+cJP/vIU1ww6AOlTGceqx1YnS7N6t8SpFIcIGVIf7
l8zdQBkrPSavC9xBw35C+dMMtIBNJs+9gKVS8tGLLfZTWSaznPwsG6xOJZDfWfordCIGSBxIwqW7
FGSVdwc4
`pragma protect end_protected
