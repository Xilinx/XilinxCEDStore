
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2023.2"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NzLmZt0/iB0aWRCqQwNeh5QRIam8BpLVxcTtL58LZxfHdgBxVfFV9cGFzr8ZvQIIinuyyjS7eJY6
bg5t5Gfu0G8fpXH3tuKOUMEY5S5MBfoD7qrVCOfsAMCccOPkjzpjwCURhJ5uKASweC45Lwe+L8hA
VARJjnJC8Qk3o/1Di5vwQW0alkUWxAJ6ogfuD70ZxM0B9wfRRXuIuEyxO/07AURXjAWp7Uwy4aH4
sTVtrsqL0qJqWzDWGi0KOTws3/Ts09ilX+oKJqhlNglJIt+J3dp56ukXlYFSCAUf2lf/j/kkqeoP
CL3anDsv7b0n8x1exXvOAqhRohgqJPYbdHK9ZA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Pg5Zv+kQ2N2XWz+wNscZIukX0JsidBSNbfye/S36fezhRR45REbbLVGxI18xJHAeGTXGh27r+2PK
9ZC8NM1l9mpc1gSZEjWdYuD97pb7MtTqdK8DyBYcWeyWVunhI14WX2ZTL9Tsyqzu16FX6lrJq+J1
6xA//WWNUqAm3B87Nm1gvoxpKF51K8Mzuh+57y491eNDrDWk3v7+I8gzKRjlmLzrpRB64oIFABsH
eWYLMVZUXOkpmlB659zFHDLea39HG5zfCzsQyY3VUmxs7pf4xhydBbvS8qIJd2Wf9sPV0LUDRhJW
otMKQyaxb/57CEgoZZ7CT4atvxBygg/2Pk/0kA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
eCvDCcpaYFOFtIL4xFaa/lot40oGQTL+oZwKLiIL5smb+j0cRvpQwCkOJoxu9ATGMl+m/yqbRlwi
2kbs2EKAB80uw22uWBMmNoOwImU9rv1YnGu88q01FzW2TRiQ1Bu1U+QNwrQ+qQC/SuuehIW4idhY
oNlKIcOKuN+nKkDjzZI=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
xY71ePua2vUzPsJano9FBU58bxzwSVni1nxQ/FQRayFfUebmOw4XxEDUN/fCq6d37uoUNak1MEkl
PtUhjrq0XLdlX3rAm193IDBrGVWByK+5CvpjS4p6P18yEXq0wCqBfah7esEL5x8lFHg+HjY09W7Y
sxuTTzQvaAGNgO11wRk49/+eIWz6H+/twIt8Vj4ZVo1NOVyRDbr47hF4FKsBrLm5U2QYxqXXsYFC
r5lG9oU2DRSlwAa/+Zzk76N6au6goxpRlFn5EO7QwYq02J7Afg3tUsX2lBkDTFkhncanfCteX414
cOC8cNPV4jND97qk1z7ou/dy1/RxaYSc63XYQJm97ONGdjx7fqNiYEN1GLwiL2+xtzM8prUk7EJ7
7zJQax9KMzVKWeXlM8NtWpVS7b/nyiWnDF94DM4Vms7ySAp3MeL4c03HKSfpPa9Lfxyt3yMcHhXs
FqM8jGe+JqX7SX+9Ffnz/TAUJ+v3UP/zouIlrT8H/Egq75ncQa8WYmmaor/UWQ9wljnalmSGM+1h
gDtSLaVdMg1EELmMWTFxsXdxDD/lRKxeBynD2yc7JoLQpXkOZW7SQyOf6lOhZOhv/7IQWQs0DtI4
3UleEl/r4EV9jPLrY5EVIidQDIweQtJATAZwLajz3RO5bIthHVKfrsQ2yy+kWjPAvRhMOHKE8RRV
GAgI0h9pdUK11G34XmbVtbkK+m1nX2+SjTX4Uegi3nowM2xcu03qs6UX3pWSUTbiy3b/7ygivOGO
Tg9bFuZckMH6rh711MKEcoVqZdg/43oKeR7yMxyHalvFpBcW+DlywGNAJAEs0zUV2aZhFn2GAXUg
SCOwunmcMG8kwveaaVPl4IPbdgjdYPmPnxa9Kk3p3TkgLFSWxeFsJWQxKxVcn1G971ogIoR74NP7
6rqtrS215B4P5cb+lNZdOyxcUvwNvC4Q0zJdhTKRXKco4LzjGEooQAtwnB82LswWIyFRk6xWic5s
lvqiQkKUIl9EvuX2Yc1axql2b4BZUCxpgtF8BXq/Us2MtGfheZeoPw5ZuG/6jdq7v7SDHRXeZjAH
WIDYWm5uCusIR0DCfm8eQngb0Y3DHCmOqbSe2zUiqem8CF4O3AxOsQS5joc+0Ohs5aJtf8uHy+fW
8KsT2xbd9d2Y+qRaLewgdNTkSr42IuLSLBaraaLxnzTNa1cY2ZBq4H/xGdH+yhqYuje8gem2v9Ns
fvbWsNN9EHwgs7kSmA47aHCnGeVyYC5h4q6njujIMxs+vImI6akKCSy6dF8asYrbZtBfIPUFacmY
OrH5JWfirTU/K8Nd9MRFfEnB8duZ0QeWWGS+LHY6xUD+0YdV6+z52mRtTI8o43uY7q/oJHDUpfci
xPdpzCe6RATdmI6NOlW11EsjKbfZvJKWZYIXQGnlyHvyZ8jctuhbuc+DdFo+nW6TNOBbtiSyAyqD
PVp0DBT39wXBsr0MxMBzu4E3bOk0Uvdpc4271nB/wdb7hnP3twhCVxIEU7J/AB4AHojnwk5rvfOI
4RYEbFvplZLXi3JS7nO3su6cOG1AjtUhk+BTahqGnpKuqpNiyDK8MiwhkcWi4yNyG+9JS/qI7mv9
OvVPtMJ7g5hXuRNsqfu+fztuxqVBqr61Ac4gMCtmTAHNkysxEhqQOHx0CtxsauORemV1gPKcQooG
cGwYlNLuWlFug9ZH1FA+TLsdm6zyS+LhT1dDEGotYlo/CcqeY+TUqnMG1H0bzQxjtoY3lIZfyqHm
ewz7ND/ngsWeTxhi2uVf83o9/JDGUiTBt+7Rf5YT+NaU7tZ1lEKNeZm8LxsUXXl/eIJvRN1UedQu
FWZthtOFAqJuxZYDjLFMvXwHRpLpmGQVpzY5ykJQk+0dnX2yv7DCRNIKjQIm315vLbpiz7xaXLTZ
q9k8eKrf44ZiMMItwCWO4ecetnioRSAoy5ALWKCCdxNgEn2TQE4jBrnL9HfsHFx4/KUnss3NDXkO
Q8mTZj99jN8XRaCuF4EYMDHm/Zgv4TrSgnulAnXgKS4uc8dbwDJUTJqr+BtY+OIZ4JXMxttkWLsk
zA7mYDH+/rZfFNEtTumrIJtX7IIn3rL3/gqLb2Y7i7Wx6kmqxoV4lxs0zc9Np0KXu+cjhE5UuFmy
xGmxAvgM1qiQq1puAmpdNuHk6lmVx7/CaLnuVnMSE/E27afma8rRWQUbYBK1T5XZhZa7C861C9Ok
OIX0qBLv5jncyStbgHbl6kXryZIAxfLDuAKp8kij5vL4i7tyHVzhi1px4kazv+ZgSeLgKon4r+K6
+GBAwr9QXFx7wywwnI3lwtKHU6gwq7CVgwFGIXOiVslFsUYcvA3APhFHoLiiYtwdBHHz6jsmp748
QCEYL7zgyqwSd8vglrZ4gAwPi9GpUVP3Bnkqrz4IEEpzPZa+eO6CniyhAMzEg788mZbCMHhno2JK
jRckTK4xoQCeTzQJaNwo/1TM9t15z4uJbrJzMEXhKsTc7zVVEfE3s5D8w3mdK+9xPwKV065ennql
0dkNSmq47LnZfGMkmf6tj7jTriPH0fmWoULPCM0MPS1OWRlyfIIdUanzK+WA09vP/8/oCQ2FLz5Z
ijWQ8dDVV2aHTCtimZrhZyzjCENW25QSg6yzDRNFkwv1iUO7BSdeKiUvDT0h+fzxi5P355MEqic2
896+W+XxAOY7xgpg7uXIxN9A8SF3dXDLEzJPUuRuvjSnptOeBbYyiG81/gK9ZdWeWZvIDyXWcnck
iz50el/o3bbJQnAmMr6gXYd7rb9SZVfmN309BalG1JvfVt3roAj+xuoKmzI/RTcwqJFydNtJNs8C
IJT2Hg/M8AuWg6hGk7SRKgZdP765BT2o2rGFQjyxK4xSCQYELesVylslL3P2KaBifEPnzBiy5csZ
hr1aXylo9OSzjiUxpezEFdyN1m1hbUKqQq5EACswCjZk/WgwFQqR7mrv9OPPzBI0cEtrtxC1YBYW
wHtkE5vh4M5RCZc7J4Mies9kot94TxTVM7w7s9YVxYlQvn/+RZNgoJCmoYpDzlsjGbgdah5yMFTN
CoFIOyG4YYFCSs4r0DBw2MocK4W/gTuxqWAA61DqXqcUBQr4R4TsarXt9juQT89Y8yl61M5wFSJS
ntQpnJWhqraU0mZ53l2HZDkZY+ryCX47Lv6FSAIxcJXSjJxHNeUEvV800SP6Aad4KJA8RpSnoTr/
b/Evsxt85oTD0cfdYPPsGMHmUNeVpEWTZ9E3JqcaT17qgMH/3o60eeu56kuQH3OMaYy3PeS+HaxU
IsiYkQXzz4rd56VnYnxCp7jF8ndLQn+tPrYX6urVIx26ud30aX5x+lMrNCK9NT3taJBLFU7IydeJ
w3voIgBswmbznJoiAl3dfXh5iAEzxh2PfdgDujleNjsnTK5Y0mX4Q/iQad5E7G9mLtb4cGG+14i8
FLIEEED+lobihSrAgpVvHofUXY8ZMLE299swUKOSnwh6Oymtde9CZOsBNPNVgrYUC8JvwScB7bGc
ohcrmlZAoi5EN4jn9zPwFr3qTUTS5m1pqqvqkXDId2jEIAHXfZbw7+MrgZBKko6vWcNNt8lXEsoG
KRitaYHCuZMM9if/Qym2Qib68+uHo4N5hhsTrmw+AdXHr4J2RzOCTQ2q42ijlFdNO60qAsXhEcbm
kmpXGLD2KEVaRV37/9wySErsR8HDLKPOkGEFYWc+9QRXjbq3+B2eWXPndco7O/ONnWkcFC4cVbgF
1KnZnYpSyV7yrHH/5PJg9e2ZBp6IxN+uvcGG2pyRJ4xVBujuLSi6MMQGd3RwmViGDUKJuoh4bzFg
SagDQ1/K1S3ftoKe0U2XO0XQxtjspARZ7NqHd8wwj9P2Wf648NSqIp5IBE3xX7NXKN6aFbxjjbbB
ujMH059UjPEF+e5oZGTx0AuARbb4pFAUWb1/S+9Kqbh9xCmshksaX9/2E0x0XzDYsNN9zKX9uWKg
Evoe2qOx3F0bSm24zw/9M1mdLUZcV4FD9lWLlGenXgike6RVva5HIph2jPp3tZxX6/bsB6MZusjo
bkYPWEsQXHXBrRiknB2VyxIxeCL4W8XtuESh9wg4KjGCt7+n4HBVikFdBeTvEY4WoFcbLQ2Q93C6
kOghif5nyTc2HWesgU+GxsxLbbJz2tguyU6+xKv8HEoYmogHkWyBreMNu9QQR6FAaEJvc0Fgp6lG
7ZiWhCrDwbYlf89JfHOWgt9WlQBx1BOOUNG1+tpspB1hx4M9Pq5AYDxDC3HQRp+LvQuDUr2rJErE
IOL8Ll21jl2Hk1bMMXN0lsdkiYMCQp60YmsM67L0taYf8CuSoaZxMv0HlRBbKqvljwVmbf3KEm8n
lmfn04+3Py5+UIIaP/euNMwrnHxBOExpBz4UG9gbbWtd4RVYtbuRkn1GZ094t5gU6zpk8/jgFS+i
bA0m+8IjqjldkXobHHKKuuR8C6vwuRC+VlCcMOAlG9HRZNjElVwzZbTOb0xJYgP/z2aRSBULuuUv
EwsbYe6P5ivm04ViVHRkFF6ZldWVupfWTFhZ+3NUxVWCKkD58UMH1dY4FX3O89TjhgUyF9yBkSN1
NYMoFrzpKDjDIComHJmfeaQ9cCG2jPv2nnYEEMyZQfxx3ecURkvSoEAq045kKUECuuyeP4QMgUFa
mp/75G1FXo9C56gWy6avehehk4soYRNlKu3S76xWq/4r5k984RuCSDkUFnVQlfG05QqJzYz9qvoP
H77wpRAtV9S0BV5FcGq1PbZl291/oSCN/kWbaUmkyXv9z1upmDTpy/EyWXQOJz1rKqM9ZpAZgpMv
Pg0hFk/h+V9DwDwZXS5JS38Jq1K2q1LCd6w7pMgUIhGNwB230IsvXTBV2PTzJq0Vzcl0TDXFoCS3
/VTvhXZT4fby6bNCVQqBOFV700c71tlPjtOWz98Shb9mr2EAKOKWX1r4qeidumuowOddzffLfajD
N9ezn1DJYNZQywP0QgmyUSWt9XCUvp7VDAcxiiKwAoOqHWzJQUPHqNfLnsgKTqntPi6WP4Ybnd3R
wAlSTyuGrlixMoKTQukGx+PD429YYadDxL1Bxh17jLlfgmMRZE2AYylVPIvv8x8tdf7Bo+Yr7hYr
OnCCi00Hk8C3Mpx6krW9kyqn1e08rdW5/vWl80kCuVhAMkVloNF/IJVSFpIaR171d6UbKMPY/MqA
bsDXt/2MJKFocMM2mkRlFs3cCRl7Fymx2AyNcnpFL73ui8CGiUgVjpzcfHuecQ/OXYCV188SZo0h
kKV/+gSSnqdFwpangGMsP7AAUf46g9OiQOPrrFaIRY3d5xRsSqMmjhsgD1iZw9AcATKD1B8uuq+V
80yWLzhekAWVCuu9Dl6imT/WZzG2v8kPHyqFh6cscMXzTA/NhCi9vyD3fEYS/Qov+f+CsDNqZJhn
Pn2bqIpKgvI34zHa1r7Cc3mx+SkrK0K8zzdzOyHC6UcxA15YhYfRzPWM4iDd30SNctBnh6swnyml
ySVdpIdlahWUaCIVarmg4ENvVcwWuWvtuMxlbUnlnbC4nFH6c/KAxmvMx0L8vA7XjNiay32R0qsn
ZJyfgSK+L4xTFwtWgowmXuLYnhdfY7lFpRUrH7g6Ao77DdMVXmFh+xBNcJxctYtHtlVFt0SodSEK
v+SL/Wxh6ghUpNjrkP0zuWhBiKGYNEtLhN+wu8aijti8MkEhE3bMBTsBzHnjfa0qjRCAz5tgTCex
vhDv9z9XvjZMc5nQOXiLUBW7xn+1NcdSWPfqnH+3S6sjEZDUDtswlALkQ4dFsvGMbK0v72K6tMqX
HZB/mGIJmTz5SZfkkThw1WSkq96j/rfvV2p9/TrI8ry1BNwfwsZJ/EqehbhNWbRRapiIdBsH1KyB
Bn6zjWOYzrD6eFXO1jx3n4Kj07xR8qcm4erCa6DhZ4q4OmjqPVE6YJjtcQLW0G/7+TFKBCjx/eLO
0UOYgPsaa46DXcfdPpKAayGn2vUwBxqvM9Bmve8XO7Ze9XkSVsEM+L31SSbr8HXh2FWpROc04nX2
RRogSV59Iqhh+0bFSq/Wd6JLXgyrWiQMt48nZlF8A1b0SBQdG2Q/n9mBNWcoBpdMLkw7GB1tfhdp
qk1d2XMLBcmZ/9NOd2Di766l55PK3Fzl1J/zQSIYfadFCPUYy1AhX8GIUXT/S5jAtT63Hhgu2OU9
vNMUDeW449Z4HabifqXVIi+uUIMBdlKw6YbtjLwj5IHedE5mUOihNOhqXqaS27tC6IqkUyiQW+xE
SxphaY3Hlx3rP1bnRpJAotDPDMvwCY5KsHnUTrIbDukHNkgAJ56xQxZQLiExBQavYW0A211GVmAg
7ae7mkY76oIKTTBrRTQfFw8FVBDGhpOm6aI1ZDspK++sybTHSnK0KezIC5fekzOgbqPDrYFGY1HV
V9OWPJWkP4Z8ks837b25xUP458kBQ9f32ygAjdjvlXJR3ZOsb2a4wyJO1oWVZO6dZ721oKGQLr+j
46tpayrPJbYb7rX24qEEGhkR8INXGPfHRV+6tWst8HBzSzR0vCDy6/WsUxulQMNnXKMzldCk7ocI
7tMv++pCVQiqHrSpy0lXaEkuFvcmcIYYYbcB/QBYBAZc7uz2JGEsv1AmyPohIFfKgcrs+3dFAaIR
rwtAOTODFkQt2lzOLhlIoFvZWoba61nxOUwt1SW5CgsYO2MDKMcJiyYdRZ0FopN8TYjZ4s8Gzk2c
Eu0lGq0L9TySluY3koCbJxsxryyAGc2EqJQuH0MmpeoLhj1y+1Sd0fr3yaYXqemSkv3zzFeFFO4+
aFR/melMtGH9wyLUOWutRfyjEjN+LwXiwNc9DqbgVfV2qd5PKsWf8Bg8m78+FmT+HG4CjUAu8Oz2
zfNppfPnlbfaquOtXJzZJQ49B50vYFr68fLJs6Rzx4jTxKf/pGza67Ui0ByFkXBsZCPedN/CYEcU
53M0BSGs+o3lEmVCMZtp0Lydah/waw/E9xABkSlw0cpVV+DG4D7XqvNIsIJ2ECniTu62KDPi5se1
Lswi9MatAV+8e7BYAi+u3qdtDIJLVT0VlDT/IQlPhet4cQC2CbwHabtx05VX8C2EmY6c9q7caR4S
Z+xZv7wFgXllPBTHuNpIiBIdGsvyCRQPN606k2TQzQgXjFY/p3wGYYKURQ8Aiih3VBMnEkXouG30
VbfXgzxXuky8Ok0ikuYx2I8hzNL6Ru/KjQqKpGpPrkz/danWwWaQhAnK73ezIK4XV+idRTUmwDPs
4E9lWgnWCygzo/dWJUQeFJRD/8RAUQfXdwXsc5dVPiqbjuzVJ6eMV1UzWe/VOVGlk5r7uOzLWtjE
rW+cGd524Qfh+sX6FXijpyrYHolwSqWLfhuvmGdJ3SSpogst/IHh30ZAN/A+qu+ilqH4QvNHSxi+
IMlo7FfnDd5YV+EDXBNIA8Jhy08qCuwO2zsgz3e6bjqwiH6OAYua3pqnZ5HdF8pwNg6UEBOfLBbB
jHD34noz3RA2XB/mnjiyDFrbxHXsxTedIkGJK20B41+879A3wDNdTiO34nFzQ4l5/Ij3E83JaceX
fDe/XA7/qcwHQm2nOc/iHpd+341stGZox5o09LotSadh47mrm0YvgRbY1EApSSIvu2f9Hq1y3eph
fpAZP60LjdllzIXfow1kAv/LalgiWZQoSCl1G5W7/o4b9F/NB0cKjZukfa9IhugeCE9hl1O4Dfi0
zO+vAChHmxQz1zeqdyQZzRurwXnhEApXie00qgqsF7Cy4ofZbkxySFXjpti+s8uXZ6U6DttTUqtR
RNxZQD1VQycoLgcwEf905zIWsjTGOQiEisNI4p3mra8q7eAmtq18ImLf/Z4tpZAEHgnkSk5eEt6I
EJQKYUchB8vMk0CTDpV7rUlHZZpkDsA3yv2m4tonKKF/d4QNyviKGRbQyfZ072aAN7SQqfFUBYII
5i+0/lyBv+8TegZQCygepQSe5fFkB/eh8Z0SxWtVPQkp1s65488fmTRQGB0ZDb8JfJ0iq7rA30hV
2ZV7NjlSEjlJCaO+So6xnxOnd5OsFbPqtFl2QfV/Lim4KCtvR/61qMsklZycuj+cfnjRAEq27hKo
pvVROZTzPQBY3PAdH3NUHq4jxqvSTFEOpPfyMWvTScpy3t86cCwuAniLb3yZGgJCrbz866aisv7l
YFtgzecGermOQMVcZFNOIxGzHUR9WeJ6jE0UXRzzyn/Z7UIjDCPVbi0a8GtCUQH6lKgj2aQnuUCf
hCkmNSRf8Hb3X14mijAb/ZFwM42fppmVRyXmBrUAIgteacHjabswHY2uIuBdfRUKwYwpRb0pah8F
K9l0B47qfvrh1ruv/PAJrWoawLc3nXiXV6Lt+FYEcqL93hw7YSvpeu1mpn5pZPZ7PPLTgggZ5peC
9FR2xw3hAunF8HV8fWuL6/eKfUXzbyYRl+BEk8DP/SWVD2o20chjaCFALD9CrY/OqTrqVqOaYQ9N
P5mFwGVxdUEoysrC7E2LqwF5qbnKWgvF1NSadCdV29Yc7HV06rIUQ1nT/dqSC2uMM572dJrs29ma
OcgiUCX1UVurWGTfzwqR8DhMrrh+2rkcMWdy8uJ8miLeYBB0aYENsiworoell+vb1u0P7h04XFr6
uoL2z9skGTHk76kB/3u6M96/fiFROmzlcniL1QX1FDuwhyD9dB8iIKxdGtXIjiIOABxXkKBFVHQJ
wOm6YP+9Jig0YNmic3nYLa3msGEiZN3aVNU0W0EuXRq+N+/oNe0figkWN+Pntun3JhL6ZtruKjC4
PYGuNsBCttKCy6UF0c2CTzEpe/kmysyN+p79wt/Ow1b71l/i1S2JVIVwJjP6ieHaFC5lshKHihXj
PMIHD/avM6tnAwMOZNBcdOIIMB8jNcqAnW8frXRw54mCgB5AjbB0/wv4RrrT6X4i1nCrmQdk+4Ng
LNpwTBOPwTN78Oy+qb9FpGOHdIvHoiXFiIgQI59V8ifzQwwPLy1W72vGUjahsQDMH0ZXsVUUvyJE
sgYMTY75T8c+JUEN9bN5slrTDvtNLGOO9JjZVFHe8qqEsywOCeewe7kbVOxE2kYZcLhqhVVHt0gJ
rimacV8gPHGxwCRcIilvb6rJaTmaeSWnH8k5K/KakG5HKm/Cb6XlDfyYCPuiomxf8Mo4767MISIC
VZvTzgTu5jYNe5a+Jhw2urA1R0w0opbmkIlde4n5P1KR4UcHwqn4qYHsTxaaSFtahIjWiFEIhNkC
Jy+gV/EEl38sr2/JJ7pQxwXkFMGn6YtElc3cSxwn3CcxmOkv4CHaRmjgwDrWD+BlDEUmen4N808S
YVRshHpCzecSLYSyoR7Nggo2GP3jPV5C7I43Wgdj2ymS+WOXI3vzknW8kdyH2RC1MrNbjxx3E3r/
gDg+wyeKtZhnNABdmDGCfZ8DCRGBs/7IaQq8MwkIJRlsDlxai2dj3xgEsxxemC1fPd71cMv9UrQe
4S3Z5wqSAAsTCY3jKk+jvJHwlu7NkSFJtElm+IROkKJgnqyn3gJwHNN8H2E6t1FlzhQvfRTH7vXR
3kuBXIIKQn4xswW/XKnj9Ct24jd4pp4wDoyRn9nF5+XXfg4Tl6S2l/BkkxuOQX0y+xX5gyQKmIwi
9odgzyXnJunfI3fPStL+HY9XXYndjaZ+i7MG2zFLZzRLQwdI9Xjs3lMoOwz7RYjlFtLBTSjM9x7Q
GNCYoqnvzwJK+6gS+p3rYXs/StX5+IlJej4uFu2Va8EgJdH5MphG3hUr1fuBF1dNhBWfENvtLY9h
RfIaMf7Baj6zqt/p39zLJOab8JTBq2UbiL3AUyMw4/7AnD4E8aj2M+Kao2pjztalTtq6mFi2+ElV
GJYv4VkrieTYJDl0irk45e4/FDnwE0ZSwNi1XdLOw1RsxACh0U16zKIg1cOJckSJAuig4j2qpX3g
AGiHN6bIWIWgi4Soz4F2OlS4b0Nfh/tx/e/w9D7zP39dx/dY5MfT3J1rbs+ifFygiPRqOZgTjlqA
k8wdj1CHxgIHGpJLM/yqkBr6uCZwFuw3PCaWemXgZ85urZjMF3Egs9TiBqLB030OhmR3a2gVWEOO
kx9CyOW+rcD+3FYCTYrzo0ytLoL3H3XWPJBx3kVUf85HZDfnNM3GNa2nynLgDFtzvNZhNcDd0qhX
STLRizF7Gkk7uYxpOBrAtu7mTatcimjdvIafpjHv8Ve0NTaJ5wdmaiQmtlXjLCRLWrkgCoScjzlK
Mh+a9Xthafxc72pADj+c2ABnc5sShLzyaR0MIU9C7SerLEkd7bDK1I2hT3KL7SQjV+66SmVPlzbV
YRHuYa8595J/6Qz0jKjW/403TVwiIMeRFAYEoO43O3n1QzjAmVsmZ1aerHLXaAo/jWLvWHoqsypl
WwFVvKEoHeH1RXDJtS0P+/zsH0rck8o0g79oOiqa+/PJsE5F4gzuOoaL3rcVm1DivxA3xJD3rpNg
k4FqZQj9l3Or0gV/7kb94Q6VOZT8I7xQpiul5eiRvCwpJBQwySuBRTVTMMWZOd6kYtaxROmULA2S
W5kkBrwbpMczmX+QOfwCYFPsngi1wH3QMdzTe0w6f+qF02l45zRJLVLh0ARwsI4nPs4IggfIEZCE
Ku+oiCebmCpUiDMeWlJorH2WR39g4JKasbattc8LUGRO+fFzc0lHgAkQtqHfX6mfmtNiYzt68p/Y
sIcXEYX1U7UNdHDTYUVnEtAH4tOzvlI3m9rxomm7HBhX806ucHuyOiehR75AGr3jpZpGXy5FcVgM
s+K+0FprNfBae/UGkJPuNTeKKJmsvd7xc4IFC+6+I2WANJehm3VNtL2sO5TPhm+sLyTTtYlUGnw2
TCmUT5LQRloqOtNcnfukxccysMw6V8B60sr/liFR1isPU/fFPALzqPTwF47Ku+dA/Y9r1bEeUTvg
TpeI9d+C1IHMwH6zVWPunYQA02Hav4jUimI8dXmRC5s1wtDnvf1m2vfOuo3U0OlnTDSjPkIAJKJ0
uzH+3P3LIB340/YmPuP9+ACl/3Iqqya82ko36ZmlZqE+Ow/2M+LJn8Ny/XiITzaGvbpNPossqLbw
Le681KxNW9+k/odrqpkL8CjUzMMeqyuTMEHistCoI3dA2/zec7hJSiS1dE68Z2kXp9is/q9kQdhT
n9rlqGRHHzc8CmJAjjJyPN3SCQqEEv9BJHCE2+6o3G61H273Pl9nOhukEVQoYHJI4jMaCbOqcP0j
3ikQomVStcyHiD4xD9Puy4od1Y4ayCosKIXYzWuIgXRLtrQGgH0tZbRSeKxYDmW6wuNCX20oQAHo
rIgjhWetsEc83Sz5QsIxFOfcVRK0f6gUxph26opVusWbKCVUDA/lbcy7pSmiJM5kE8nV81y+LAZS
6nJytHrpvFJgnl3KIeHG+MVOnow6N8ANYjW50efzgvrdIQUHhf69ghjKse+PBlAxopliML+J/kWS
akQS9SrG2YA15E098SGUeOfoYndLQ7UHOYk452IQ2ZLAEjCH53hKgWllk9B1ZWdsGM6HCGYdA2vB
+vDq0By4E7lWxNuoYLoT42jCe1nyFvwEP92cKS14JjXftRHCA5Z/ZHnadI55Ws5V0Azsrt6f4kBX
4hGdMnoqixDsCu0giKZlwofO94a6+vg2KwOLpS3qxM0Y/dWcDb149zusn2lMb2oE+y6pVd09dTh9
Eib6mLHXo9xIX7lWcjqwiOLoSKjITCfd6YpB6SgStr06TyrnK9VqqYnEdu8K0DDZ6EwgU5JNuasf
NKSlwIuOPFyQdXDHZJEGefMU1XYUUZzSLkadInV10pJtdg4wArNgoxCbUQls+ShLciswDcyCo+6m
lNgVXkuiugiL0vjyufpaiIVBbpz67l0G8TKXlvswXMdW57VWFzL1QEn/xXDAovl/i3bSmU6RnTcl
L11QP+AsuxcyHnq38eRQiTKV9eMn1k+mneEOC1kqoxYzLTM8FOD5oCZryjyxRZ56F3jCtp51MTAh
itxdTs8me406j1oVWImtWUOQ5nzz1UzHQzaWMj9GaL5Fm4kgCxpSH1RS6ThzJ5P50dnKzscS3Hu7
rDrD0UA4fuAgsycdwc8XEeHxGFqHm387aOjIKGl8mz7wV930l02F9fNLci+PB9BR2zDsb2cbTnZI
x8lQPI6Jlpz1kVp2MdQZBiO3ZEoBIbwgi788ujpTQNnlW0MMfhWErCf46VN3BKHqaHG+0LlzYS/U
tvPviI8x0rdIMAy7sBZcGUXAIpwMXd1ZDD8ipEMKIN+w87tvo3y0N6yi0LDhGt1UFu3LGH02D27W
gHrcwnCVZD8JJlMyRRQ0h0EgNzm0RNMS38XMO+eCLaEJZNUOBgPpUaE4B6cgo0DTu64zmqR4rBaL
+o9LlaM8XgYVx1vB7HpJOX7d//QlBc6ZLqG8tzE0GzEo2kHwdXIF64u2kVszWtsao0EqUIzaLHrv
7hoV/AIe8y2MN2btjhWpncEIbM+B8fE+PCrxMaKGvidxYZOJkVWFvORB0iNq4362a0gst6Qn0peI
oq03mg3ohe+v0eCsCQvGtPgW3stIvup73xzd1rP2fsYG8pOY3gUWpET1Kbvx0fsl8eykufPEcPSO
bsR0so4Er716zrmzd5G6+QNQjXvInKuD/sTiP8612vpudCS3edR7LFhh24c9qiE7qaigylm2wbJj
/d5ZHudIo2XbIV73BkryFczAU0LotWpOEiNc347XsLSEh4IQQNNLSGcl0+z5H02cV4wqAr+zvopi
ikvXS5mQx5eJi1MzmtDxsfZDIJpyDi/zFWHtl6/3bZPlTvoEqpg+iARO0dOi6ePxriDH/DY5CRXA
XkZvJHKhJPLQKfxwogsZD6XC1wMXGMAls3QldyY5MIKK7f7J7BaO0CRCGid6mqknT+/DfHXjPHI9
+Pek0isiP9XF2quOS9VguH8l61IHuw9U2NN6XszbWrzvI4iMs/iVQEIJiW2OrgutiB/JhYnFn9G6
CpTqhjO3s8yWlnMAGJAY2Rm+3OIWEcsQfcVdj3UATsuqtHDmEnbPyxhZ8BSFpPthXZ+Rwql2/TN7
3wrym5jmVwwgpMw87Joe8P6TWrNYbEwekn+xoqPUt0ILDRTKaIHOJ0BqteHNL3OoVurH3be2HZoA
t01u5EflUxYdvcOTNy1VjiPMXRDmf9rp2tJj6zNeeyY2DJqjuJzD32EGKX+U8+2f+vg5GUlwtEi8
XskN2Shub26Huoi73X2o8xXtTqbEpbpTkjy2sAgAnd4fkOohfyjctzSpXDtcndqMGgewDRLui1O8
DRUNPRD6HSWtzk9MDAqKwMSpzj8mN3+6zi5GClnj+aYm3PXRIOxmOY+d4ZMNpN9nW/OwYzJgbis+
ckisnZxErS8CiDpvSll93lF981VjZ/LG+c9JpyNNkjj0D2FcLV9jablaPjdO+/RYS/UJHGWAa0ZT
iZTqGD9NCci+VJyGmlUJ0k2R5aL6mTipLZ4FhArMoC+if3+kVHD3PN+juaHh50lq9o+wQi0pQuOH
/0UjLaBG2h8b+vISs+B/fso4dAR0/rLmhtz4i8MJ+npvcSTIyy0poLS40rdZSr8RbI+/RNDRypir
GBeHijVli0ZxAjjqdxGIkLPAFRImd4lMFz6omi3aXp0LssVCh7XissITq2Tvu7LBoHBWO3M/u/RI
81M2oqzWKTSKHSHW5f1gQc6tyAIMcEBBLLcEnKGj3KcPbQTNNyzuZ8qf0RKY5adVdSGDmg8W1EBJ
i2hCpV3VGtIfATw8kZbRrQ/p2v/g86tlpA2a8w304Ax7s7MeTJMekkCwIi0EPGijkFIB7YMU6KzA
xltJRy+0PsBgL/HQBJ1aovtYsV5WMWuhxe1GqM+rLxqfPGFJIUKxBEiGzm/FyQkzuFxeiq+YlBy9
tPv6pcDWy11LnrsHhoR39DXV579CqDdBUr/jcwMVClr1poAczlbcv0pzSTIvdrpcGFeDAIUnwymX
TdHIG9o8DnhJDUOVhKG/yLTXy4SKAmjZLIeTiEZCfW08HlO2x4hpO+s+VfQUWuVAlqlqxOlh3q6R
DhTw6Cx9bxxIvU7QvDUNF00353qWeErn/QH5saTtpFS7V2TB1iocwBmBFPiLHBQLhTdmN/OG6qU0
Rbyfagujw0JCw4e7IJAcGEGigaC4+6buOdEoueSSh70ecEFZ+VZuIX0qLJGwiFTtQ8E9y83eZ5/g
Nd4E2MXGycz2EQ4MMBWwJ3HrMrdBYVIey6RmOQP2PWh7WxChahvkG4WoW7VS+22+pPg4MLpTOPoy
AjQ+yXH5MIrcWUK0iFdyLEFzATt3J75ykp9f1D8eqmL2JPyAnKnk2UJeE1i8waRQ2GdfC1E7O2H2
GfT2wAsJO/+0XsR4gPROCab1O+OqAzjuQI8dFCXEK6u8Pbv1SBf/9Gcjz/tZPNcZ8K3NB8FGUVzc
gTX+8LEuBJMVNPuhUYFajIMnVrDBqdO6OvcCCJ9xkGWxnxUmvbXMVI5Z/+YUBEHhv/+d4EF3oUD8
j4zdfo+cdYVKq+oZXkFaCtjYqIzjH8MufBhu2s/q6GwfViTjV9JYZYNvNjY2wMkbQN/nIaaQkTZR
/cLr4Km/5ohg9ILLpsKfyHBYJnNHEfkxflDdT/M35lPMhuIzXUdB14EbLuLzacTeL1RFfevvMUT0
rg9JfEOPA0riocSu3bNQjkIJbkBMY84c9frr7Hr0HfZpibErVyKdAUnDYSqIZ3ZjVBVlqtTJPSlt
pBXc+arH9qmLyTU8T890oiHmSzLuGaLzlPFX7XmFMWjfbeExWnpUN1IBuwbUKaiyKBQUbuXVSB7B
MF7Jpy7EIIpdLW4vWM3gpTOyEnxUc4G7pkIl17/wCnXqyjh1Ov6UMqpPX0WrTtW7mKpdRen3IRXh
uwFB2P0CNRV4taMc9cCcnK+pccDLOhbzbPyw9Fu2fIRg7XEybz6V2yYjXYiDTseeDkGP64VqOW3Y
TnA8Op0pFeOz69r5DF+RtBc2nEfWeMksB5L5j4FA9fZHBp4ilX0Nn7izSGN8NOUfKnDNqjWcsGd9
35k6wfrP09Skxnskq8TkZBj0P4wHiZLb3b8e8Fc8Wg+Vi+EB1CDVPuPvumb3KCEnOxJsZ1bIeqgV
dQDik09JMKYh8eXNMybJJJ/NIDyAhpUzkpeVSfpakrB8EmYlkL0OBF7PE/yL+YDScR0X2K2y6dM1
mT/fD9LZ0nCH+1zPnnKq8ecacTOM4ROQh3qMdJ9GRU8d9L6OAG2ww3Edo+7pa3T9YPc0BTrSi9El
0nwQl7VhhdEEK7AB8O48Rmvh5dMKwMhFwQTqLecTlKodRQPQ0tY5cikmC1+12+l/cLKEZ9/jD9HX
9cq56mTy910O1y3c/E6oShyL57x39IeLC9cahX6X/9CfIeMU2YOer9CDN24j61afnfyYaXBanYX5
gfatGrzHRvkNM5VvzeZ7YUQquZPfvr040Ylc+40vQ/g+b1P+GnFaFJk0XpD1XW50HB2FmkkpiBbL
uFxynsnhKoJ9K1/OI10LRueyehvpfQyNVJK6pFMn/XEKFfoFPkxCoov860C3u4M/2tRQGnRk2Cb8
SqMRw3Vxr7a9AnSDgW6PrfTVU5NG+DGYXOO5dL1fG/Q7//zn6FI+JzVZKv85hdU9hl7QceyfJMI0
XP3BsEsoEzY7Z5TOgT3qmPb5/cLRAZUyDjVle/BFhPFCnykVkMkqxbnViTAI8qHfOs8taDe3yr7c
RRK5aPtEctIqg6atVg3R0ABRQXil4q+yX+JPx0qXSqieDyTZ7rxL9Lswgw2nKYUeWaJeiaYhnxdM
9Jf53cquw1lwswTemWuTj7v1+x5mmLqIz1zkkggf1kDE7NtpR3xD9DeCohkI/0NpBAPLIy9skJmt
XDJMrlsfSvQvCBjVjefQCizrbs4dvNsxIH1i6/ggeRlugZJS3XniqJKq/RsfnBhc4toFVDMqIiVK
chTYrlr3S0BeLlvZRl50XYJ0ibFzjqExPqbZvraqCPnHbR2j/7oXWGT12KQzv195ICc9QTNV/iTC
vEaLgyMXPSLYhZ5CEfmSLk4iISaMe/RoD6h6e/192zDRKs67R4IFXLBZvTlu92qSa1eBhXzkdjub
BizSDbY3r5dmrDYtB6yulyrsOlWlrW5mQyT16oHufV2RwdTTsWHkENjGM+mtauy9HIGjnvBgHphp
wwPYVvwZV3IDoNNsCib06mbRX0wTwJL/XUMB8x4lHbHmb1VZ+UgyjJk4Og0ejXPs/bsR8uqGznFS
BcrlvtYmM/EKJnxf6X02w836uwVxL7CMSszWJNX+wL78/6qglXw/NCv1/P7u6TPY7Ik7t9cD2CxI
DQ8n1AYkwWM+IN88YVpPRLZO6g1JZREUAZdUYaUQ0VFmuyLxsQ7L+n3K1My94+3FM25r6g3OG+VW
7FfmbBlKkhO63Oo3Hx2PAWGAWuCJ+/OJUpI0OhiJdR5y40w8ePB9LhP46feEwa7a88xgnb6Ozl34
SfON4XxcUIUfVso6bZ7Kf8jTFSNZz0z/OijAxTI0YpWlZOpC6AWTsuVf/ES07210hYm9IJ0v47FI
qBoI6qMNDKO2QwZ6xfQjyhJrPgtCnRv5c22CnOiFRUnthJvcEsGsOzxyCfN8WtVU3twOeDKi+GDB
F+VJYyEXhKSKDh3Tbtct1/TcYmAt2pKzWyZAGgR56rZUh/vzm+BYRW+Rz8I7gScNgymwYffXcBfO
L2zjF+U6rVCajq4PxPaM7uJ9w7CzpACdF9Wp7Tl5AosXF8eNbHw0QPZbJgkPA2/ydPk9IZJfzaMy
4mE42xzRkmQmgh0bwbZ31sEAb9l1XFWxMcRHEOHNwR9sL2vKISofrGESSOBtgNz6dsGputlqCom5
IzX4gFrV5ylm6zsZSeMPaT7OY7ayHX8J45ooUCht818aBFnUAT+dN3eTXUZiTeMHsUK1AED64CT3
M6WOto9BzEUnESquJVENLOYY8uX3ie+Psgx2Y0XhLN5/1YaOWKd81cE6zZFfBqVoDHFzMEZSlNnl
mtZO1JLmcoOZ9JcJnfRI7B2/wXJizjV5/ahglxjphyj2NAIq/euhQyTXzMmlz6jqNopjJQFfnDol
adoaglQW1UHXHzXKOdypdRDbuucLxflVFCKQvgA4zH4Ps4/06ArPi+zd5yVO0PXK0G0+LIsKq7dW
X/qk2whwWm9b8tYXxyClaYllEyn9FRKkMZT9KVZBpmMJoU0Jxaljcuv2gQ44uwwnTYU367Q2oO5v
epNyvM3kcq7L8xShTTYGUjnQeijWKn6mjK6+xWk6TigBkiIlv26hJOXnmrbrm6YEoBOxz5lZD5vf
It5Wc4FmUGmg3/ltt8VxRl5Or61fLvnJJ5El1ucDt+1aKgREXCEyPdmXih+K+dDDk06bCTCUyy9/
mYdl2x5NqEBdrY/NYlcpQaoBbM1OqMWiqVFxt60zo3klkg5wPW7+i9pmJS/zajYP0fJcNgxSewZH
P7TkXbICc4z6kW2bkEw0lXWWtzrsgswbl78peT9+2Gb8MxQZQxqnACL3ygNv7NKPa9DCDFgjXyPX
QmAIwDCKWtZK02gyGhlCHY7l215dPTFZY6Js749DmrBHXSOK3iDjRvJiJTrbskJZh3JpbyXfarY+
i1yH+ssoweDrhrvZ/Rk1znU7QdswuDoxOYy7zgQXb7XH7c32kJPPr+hJ+T/aIUxyr74nwy5m4nZK
G+ZWULSYbgxc47amR5Oz9Rc+Kud1kjmRVLIeUsajn6zizszm1bybLNJG9IlVLqRk9403t2w9i9Co
Hrg8ROxsU2IKk4QclNnY/nYTFaaTebcmCFFWaRAqj/BNQ/0UMSYTmuTik8iHBMo6X941lOeyfgH4
Yqsxt58G440NrKMU8uAIrei2v1NNxyoDphpJN71ufD4cBJglPD++2mdqpMH+aJ7NA8YtgpVrikNA
jiF9I9RePqemZY0hpWuBU2sEI5kZTDYP1M9Bjmb//d9glwb6/JIqd72MqUg5KaIFoL6HwXxmQcgb
009ahu6wADbDdVbCQhVwVJXF87TnXLK9RLDRTe9WbODBI4lGaG2KW4e9MsAnmsXcMzOONlZtejT1
Av3I3UEybItBtI8hRUgxc/Byk7C9o0qHkrfTskjHtcxLjxPOM+2jkYCReiIlMB0t9rUsdtfj7Ea6
ZlArTcE16oI4188oWjoeCbZ/NXSTi+A/TC/Ewe1x3MUBJm8lcM1C3y0muNKfzrX5Cbx4HweP/Qst
dszNvrec/FuZAlu+fJx3NtGxBygxHE86GiP9qU9v29y3YbFwdqXBvYyyii3ASwGn2TNwLQFKSGsS
24KHMGOCH5JPRviznQJLOLcmf7zE/qt604oxr/kOUMo6uzsswfdSMfa7/fB7fdVizGZEq5k+M5nH
aenAJA/n0m5hjWaXD+MXuV/PGVacyQgwbKqvkLBBqkxyTriSS7mCj0XAkLJV2OaKEGC8f677qcxO
JYq/rAIY97TKO6LMg6qP3AgjmmbK4usxNGYmonw1SnjD2j9Wu7pWcv6tDUXlegS3922Qvvk2KiOA
JmtSL135CMvdK03uISChvAfr5HelDppMh3VIDsLw0HKAKx0eMfqsL2Kq6fAJ0v0OXp4Kc24rPzSa
d9QzFDyfK97UzFVVejiwDZZSJrM+F7UmozfTtcdohtsdVmKcd1hAExje0hp4Cz4GfuxRFTNiV16F
fHORHsjL9vkchUr2F4s8bsYiVM+9Llr5wrPcFR2RHq4KnMN+ZBX6DwOGVIoLnp050poPcfC9wIGE
635ExYC1EAYH04WY0arXIHAL4JuPY9A55xGA9Sip+/gF1DJC0ilizDuHSwhCDenl2ZtHSLsRhwpe
KD96pLj9pLhdrJU29HXg0Vc+hWAxZ0ZAk9zUjPihcugMbA33+QU3/e1qIvJP6AqVouT2EaoZ3Zwv
TPgtiu9ckNN/4Aa9FoULdZOUZ531d4lcZ6A1rGG8y84ndbhcxVz/1WzdoHeE3HB+A/AfM7CD6bD8
NT3NFAEy60hB4Ek7nIc8zoKK5NYn8B4d2aCaKHAhXoED1nR6el8rbBFMDCfsv7wNbN3BTgCLvmWn
v8oVpBpHjc6HXeZLrxpW5AJ+nOuZ5oqFGFC043WlSQPBuUKeQcJ/M4gFPnTtL5JwFH5idozxQa6L
rD2riL+XaaOOv6cLAGnimox798DjiXko95VlhFo4tDKrJ4m4iumQQzSzGhEaAHhvlCx6KvjyzShb
47DWr8cVPEkqVGehZ/oobC7FfME2/6Iiih2OaMnlICu2kkFHu2Zc80mH4D3F5w3LkzEV5I5p1zo4
/Unuool1vw0EaCYEXUVp3FaYPzMIKYbVotMpCv9bm8D4kQcNZ4j/SUlPGcBG/3GaR1sUZaRsislH
spqc1BAenxlasgcR53NY7g8T1KMGQ/sTu4MjJiPD04zi0CExmk1ryWT71cFzqfFR2SvgD3+yBeQH
wh4Zx86HBa2UaFWiqgcNlfVGIU9NC8QJV6m8nOsz0rC0g6bgJqZA2vq8KbyrqaKLUtFH+BDaPUQt
MnDC6DUSH9frXsBMGoeFWh5rkw3N/+8+Jk95dl/jJH/kQcewmRDRJumvZXAmujFKesacmZGyPCut
UTmn28lDlkvg/6cSHdKIhIDIGlzZI+lRQoR62UeSm4TQ4hUrGjNv6iy6JCyvSKz/xs/r85cfLvC4
QbF3HAZxZWJHM6FGzkXqkeCEyAjYt8YvBfS9dAX14dwNZakX2FtA6Mq1/wtIvmhhi7wBWUy1bZ0K
CtLY/tWNcH1cZUIUB8vBHVtI3ZnS6HKKwtnhk0ywT2Ol7p8xuTqlPNT1yurrZjeMkFA1C9xVDGlx
IeDEioZcO5C8BLxxeJOXf7A0jbd0zF1zjwtGYBgd1PS2B2givORiIkHys0C7nHPwUIRPe6XXkA9U
FijZyMdfMg9kQCP0rrlSeUwaWS+XLTXrn69vf9sZLDy26H06tMcJFCRBUUb/JBkS2BBiOXyMoLNS
M+t7JES0do46/q1Ayoa3al6eGfa9RzC0qki1kfhlb6oFnrhTSpN1XCGodwU9QpPCUlENuAU4vpKo
m4b1XPF7fBfIVw4h6ZdEybKvGCfAjW10PH/Erweh79SGhNTMNiREjjPDtQ7+b0krWL3p4Js5N9Gc
ofVbYjsGGqsW9o6cmi095FNr0oJejNLtwGXrXoBjo13gQcbEq1g+EJvY9Mo3Q1Auv6XspsVW0GVp
D+t8i283LuqrgwNUTSBIE0V5PnJszTjVU9N6+7ka6tULSvG6fz2ASJT1wPf8jd+dUAMg8XylShDN
ygkLiyNBrETt2wLceZWkOHWThqvGlcvKcJqRczHvlOeNOkx574NogrgaVfb27ooTAo7V1o15+cMP
pETBS/U5qpj8q7Z40Y+gw6KIyL/QBhVXZsktPaLHiWSvbGE8Ng7vpTbrF6mX9KWqhjGECmdS9CdY
plgnOBT+aItuTxSfYR7DOgASRfywL1Xz7++Fg5hYESJeM3/T+dlhJXV/s+nUJcikr83J377qtN3h
v0MisqTIckZCPgn2MgjHMjZopfOZlWRX6c70E2Yh16nOUf7BH3ue798lU3oIILQUf5mcNytjQGIg
10zdAIP7bQcduE/57/i7hp68oiTEGcuOtQdJ9qMUfjhJkz1c7eS5XA5M9cokGfsc30rGnL1YLeJa
vPUd+omuPyKB65wxE1QohbyiGwAzH0IbI5Cl7DnR8Lw+65s/iZpqqGbpY1veIt9fOo8vfeg0TNiv
uCKdVT3UamCzJplNTti2qlHFPXR/CrMuIvKw6c7Xco5RM7OKrGaIlrQnZxsYNbyLDPFUEW5xf8FY
KIeYeV9s4MTOM0J5r0s1sYYDD4GxNigkZ4olqXKDMKpwYIqnJiLURgj+/1XC5GpmH6w8p2Oc8Yjt
RpWAmtXtbrS/geXC16w3tDfPeHaVZANvUUgseAwKzseiJ2SorFGTQh67cl6rJs4x0vVNxEVP+0A5
ou5m4xVMivdMgb+a4o+tuyp5hpccje1tHuTk5dxREPcx8dSiOA2vIN25O8T/zQ6SuFPW2+Ch42pJ
kPcSlJ8GPMEXXl0PG4mnCS6DmM0JwKC7ZEaysJcrBqUqj/RoJMaEi5m2DJYhZH24S5ZwjOfFpcXh
RjYhXAwYjyY8+4S2nMA7Yx/xVNW+LgLetjyAWaSsrwCxBWJ0p4NjpnKo9plrKo1BwNqpIu+sW4SE
wHOEcafQfvuXNn9SBaM/Ik8MMLWC98mGJ5z8M5/36J58Matr8PbNfEMTG8lCMkjksSpAmJJoFajI
g1o7RZ0EXFyFp4M+vFpuCRNQBDdeacWNPiMGWFLWt1zERubFycqasD8rAU6bjl0Bk1T4TFoPUIC5
fgmnmaZ2Wikh80tEYCOencHi/KFDtymhQEX70lfSSg2F5eqYGSbCWDRhDLO3n/LopLk0gLgfowD3
rEr74TotqVIiOrGYtFEc4oOShYTyW/0gUf9nha1no7O846gzQT2SEUhRtbk+jc9W4jwvNSDkky1S
TQ21vwUiXfeVeOZIW9ORQypXFfs1QsDk2zLTHjWtOXS73Lr4MPtHnk0coeEWrQb3SP/n8jwwmpeF
YPVYbRGbO8BTlwGPTgf+SswK77rPRsMG5uh0zlFliLbwQpf8ZcMLv43VYXWm6EDs2vfNmHMDORBK
9OdbjLFBaEdo6gvxEU/GeTXbyfePMWm/U4s1OhxZIsxstTJSUhTVGWDRFBsAS6OOsErz146WJtnK
1nbKstjGi9glZ9OsmEfZil+lG7FSfHbsJuXUNISHk7S+m9Fz/SY7TNVvoDzkVgUIyxEybcS6lbZp
knxxQn5yckufQQfLn7Q6c+UnrdIkTJNrLcdW/TGpBNCPv3HeV32sSyKk+osp4A9mFPv620Lvc8iz
stXn/FOxRD8Imyk+Euw7Y5qnS36o2u9+Zu7rYEGhDB2QeGE/JLWTCBumHY2sxYb3UPl1lpzMOXQZ
QCbCh+P74nvMJYU/6IV2XoYou0YMVXjjGBpZ8wzlhiJ1ugbJjT5qNc+wHLZG+fDWmypPwBg6HSdr
fxIvFeNdLxl0dekXL+gBZp99j8nsBzdj+bsvMCNlyEgp0Vuo6hx9C6lFv4f9tyrlatK08/xI9QuY
F5V9apAMsmCYvs00Nkawak5P8zS+notvKG5uy+gHZ0zsAVOWnb+fBeOSCvJKd7tjAMavkim50n1j
1iMLPGfMTvC92bDI3JF+QvV27dY7sGqoCsV8XlzhctBRzGVf3cd+bav58OecWuXHHfXf9g0u4onI
Y0Pl1qZWvsWLqRz/YOYzt0iFltawxJ9VIc8O/7NNtmfqJr/EfIwBkblJNeX/tIAd9fVoterWc3pj
UGwX24PSoUx5oBts/Cgpyaggwi7v8tuuhHlOaX1Z5zYRgP+fMsJ4hcG0LkDuo1TDZwp4XBHqtgXd
gkfTUFKpqyKACHVGe/uZuui1F1hRWrHYpX6ODPdWzvtzPnDztkcoUrjFAd5fhsTgKP3IqOYCxo+c
H/k3bcTv/Af+RbMo7PGzd3tH43HBWkZbWhlXBKXaDV1ZGX8ATKMXEIoHxkaXIFISPCOnL/su1YBl
sqp9x0jZK4jy3278hqC0DpVQ8BSrdSI/tSwrl92fQgFA7W/kB1UXfedkmXNBHeToiZACjEnjiBtE
ZmMRQmX/AMdgD02GaoH+Ryq2Vt1k9Y/Gzp8vpWjB9iLvkGXc+vCWTT5GmzAml99ZXveoM84qhH4W
S7IIY4zm8XbnHdocUJDgasdHG6B/GbIi3h7Bop9htc9UP8cqEwvwR93mDnAqXW+7e4yuLovh7ALV
EmPgFUvQAI3gnHJGIlCDlrQmgYTahbD2BsZ+Y7tAgEruLzV322CEQhDag4fGuNciI7mnmy+tGymv
QQ+7bsafWMcPRS3qSWmHZWA+A5rl+MAixCY2eb9Md6JfRadVBG+fKi3sKWe/PNTsCZDjPnYwVkiT
Ux+knWhKLwkAj0RYG6o3H9+T0FTe9q951Y8GkAuVpcPqr5Frh9BzLrYp0kh2wg4oo4TX+/Cwn3fo
2ZNBtr5qRSOZI5QgVBNX+w8xNZcbYMrzMHoYiWFVm4TUmRJ/3lCWFFYdxkhPL8HqRpM0B4FNOCsb
mc46icWqcWHDeqGbe39nWHd4ySi1d0Z1wYDVO8I4+DGnvMCRtrsD0gVOb7hgBeRL6w2omjMW1F0h
BXG83AsrwoRx7M5it0opZvky8qXR4LtmU3Vc0pftXFlylXlJ8dB6+P/iP9MYSmHfU5l+oXllKV2y
2N4j9ByFp7X465jC8nYQiEm1rJ87B7w5WGne2NbAT7nZsmz+faa/diMQKaGPKmVdX1K4BU3wXFNO
2vvpPFo3536F2pmFRQacjbZTvdHsVSu24aLfV37rOJjw06WwrbkE3pu8hyK1c/51HbqGm8XDDlCR
Rfefw98iu1AoMtQNhj/C9pxLgxgcVeDvQqu5MhG3S60R8EKYHKqNb/i8d7Zeu54Itc43K5EHccJt
VOIoC0WUVqce3t/NxK+yX0xiVzWTYOhm4HpYE9UMyu3baWGoyE6vje1P8ZLpLuLXH9bDPk2RW75f
Ll2uVsRHu2AUdb7j6SOAFnvW7sDiI+5CZ+DEy8+UiThhnsIqTdu52QqHCmByOJnIqKvRouD3of8C
xWGsPAhPKKevLISK5OUXR2znWR2H3TwoucQ46sUiqv1Qz/JI9C9vPsTI4+qepwPFijLadtxT+Lm5
mNflFRhzlCDImrV8Ml4vnub+y2z/+o1lp4IbkZ1iCPUUxgOmYXnHH0ic2byYSPEGqVeADUnSPdcP
twgACpgPFGMLCZPRWqgbBif8BGGCAxY5qbfiLb04+WevQ6DrcPBG7V3an9pouFc5opbMHvt1EMTP
1OYytuMvvggI0+x8T0Rr5zF3+C0ISIH9RkQP3T2XaKZ3TOtU7KXwWal+jOcSsSelbao4vGdMEF69
RZotcbRxwywC6w5TvjuxJDeCNNcHleFZO61QFVgwNSKCnUXyp5/hGw9KmpIc5HGiXR6+90Hsyyam
M7hOG2SZuMPR8h1qe493mvfeRnp+Ya3Pnow4rWgjZ2KBcYC0B+bj+dy0zA0NXVIF4RCM7pnl0m7P
5e5FaobrHuDoWNRfwaxM2COOG5g4+Q0zCCcsay4/4kJGr8lq3JT47TXwRmup74Qop0GlhC7dUrIa
PstIWHzJ5stx/DCoB672MgBCfbJxSzRwf8jye1avbe2Y7J5Igb4JtVC5I/OuavJMaC1LlUE4nv18
2EYOpq4o25Fn1qtIaeC1BE8obeMlmU/XnXNfkPCxxkvAiCpc9UY6d03GU/HhzysSBVmHklJ44qhO
25OnA0+OpNLcgTW72kfp4KGIeyWlmyDV1htIu+5IpK13hVt5ZZhhbHg2CwZnbksJVVbuHTEews/H
/r7mvje7pJnd1c2yApIuq97VvEnj4cUWpaEhUEQv9z6MkgvMTUFW2JMSnoiL1kZ+3UzpUWH8iduE
oud+jJRIMt/llaFUrVP5ilC1BGki2PzuIOVDMju98WoRU/Z6BYNwcppoNicvJ5EnQ5V8qGl1+f5M
IMd0NJmiuH6Ui+AMRO0KJfuXFgUBOhMMRFEwV4SJfGCPMUyRcSrkakncoUbXKm8AxJoW7gYjKuMu
A8zuqDQonUSX2CfjqIGQa48c43fhTLU2DQD0Wwbi36ROae0El5ElLVC2O0D8NhX4x9qxnpFC6W/p
SWMz4I8ik82M0Zy292flpnfeL8D2rO9YnwtiieC8rWJPAy7ffJfwsxPsHYQgITUhj1GK781zZt13
TbaEYZtcqbWiUwrARriCRgoboxGhw9XhSDzS9AhpsE/kWQpUJE7r3Xsv97Dx4hj4525EVAzqab+R
53asYbFa/QejdejM8CIbPUGVIFyWmnULHGxYHiHuvd92zvr0uh9vsXlLATUgpnLADQSApzqAwT4O
lVk6axRSFhyRogkZoSJzsp13zfhmilRJoIibHV8KP/ivXL5WoeYD212LsSh6FTmGNMEdUi+FQUFD
qYy9bpG4seBhyNg7cDPPwvLivkgb8Xb9UFFj+1MzRnK3mZ+ofN7r593C/MCdqb8Ji5W0SJKaePBU
lkNiGzv1AKMrEN4NC9BJ1aUcpK1h5Kw9i2p/F/9vbBCdTLytJIL/gq8RvUc41qNFG60z9aH4SsS6
6VkjxBr/r/EwC/9G5HZmFH0O9xDdectLjm+3thWKYfeWJkq2KH29rQY8Qq8c/CqKtxY+GYaglcUh
805jA4T5ExwshhAb0EWYlrucN6+4R8KG7rf7zV6GFstQoUNB8iD4UlikfAmbmUzn/EZimRaUAlVg
ns3KM59VMyPgVbBq15AKTM2xXoWYdzbPkwyIUgWEGyVWqWK/dHAFdD3BHOtcZg1nb119vSZpOTWl
M3v+v7ke+04whtGhynVacWLceag5fu+JwhgOLnyObF1dZCKsAtpfecvKVtKVkQUrKhTcs8XYWBzU
IVZIdqnj2n45UrIAbS4vlAOBtqFZN55S+Oxs1G0Jm/ogDAAAJqtABlR+Bxk3vpb696Hq7TuTb8KT
2sKqo4eq2BUKx//POCS6o6ZmfQVYS5saGgvMFu7aHo6ES9jQ9cCXQoSEr4K1eZiZO+PZ9LhVpYFY
wCK8d1WdwY+NJUL1bJXNzCyrh6D+RtPQYcT7eeEnsjY5FtAkG4ZtboRPYmuc960pZ9ynZXblBjk3
6dymCDybC4coKfnG+IZ4FFY34qM9EaAh7wvjA3F0k0A2hmvnk4Z0uA96VLe7OxQyzXZx03x4VKfh
Pg1x2vy7cNY0en9MmjFTq0q2ZkKLLB9/VrRpYbhJHgossTPxxcfkIltx43t34EdixayHv7drxvdh
OoohQpGMfyOLVStUHe5k43lOhTStqHB6wjl+NbTUbjy1G7rdNfz1WvYpi5/OT8oqUF2rjZNKZJZT
N2Jt9jDrteqYMFAwgTR85IA7ZNFull0qeyYgzrgHAAutEWhvL5AtABxxuwoGV4Z2lz3cxngZjSMK
CMDkl1l9vZsAj8MDwrIaOi9Gh/74ZdpHtT7dqB3SWP2Jxc31kWmMMHutj6D2RVn441wzrvv1xqCI
NNtTbWR7nEpcwsrJGcEUThZw0jYEGSRM9xWlK9LC7N9IqXDmtOTFcX1z07RGT+XjRUggs2fMVCHd
T1157HAGu58ZsHt6+du5hL5H2acP54aFe1D+4yiTN7uO8Ns0Y/ZLGLkbKz9kJlN6w9PHo1pwyeMO
LDbhdbakoFskpL44a+A75Qd47/AiPh2h2GDOXju29LRrXXFTC0Gq6NCSidYjKNUoAuicnQeMnArl
tZcegIyz+HFcx3W4RJHeNRq1rb0fsnEHIOXYS/GFS3Z0npp3xjZKD4JX9iXSJhavTY14OPhCimEx
IOXgEMSPAX96tUz4HM5MRO/ff8CZD/7vjo3c1bNyf20so5qSTwx6IOC1Bvy04GrUR939tsPxnAvu
WofMQbkQowhP+vPpORKdRiTflteMiinWHX5E2okcGsNZ2+WYU18Lk/8M+p5FV+PRHps8wz5cm4k6
lDA6VXo8T2msk4UCltVVf2pSirYWyPQlQCsnKu2LQPdg/YNbDG+OiQ8Dc5iwvt5hgyY890bQO4GE
+K1oO9Pln6t9BWOJwl7InyXII6Ni7AOtwSwSsdE3AS1VM4T46hzJdtTLpPNrdJ3PntcNOzZLRfGa
3BbL6s/5siMclUGE2MdV6g7K3YtkJZdW74ELtRonIj40ar8SaVQyOPFiBkv9Eu3kgPpTP5ejuvaZ
P+QO1ZO2obq5IJqGpiOrUai69jtBQ6B+AcgBFdZ79A47Ccl9Kbhvau2QV56Gfgx8TtPUZHnyj46a
Us0t//cWtg3ygiehXqTTzB80zefHR6Bs1gPUmJi/+YtLsc3w2BHRXuMwGDn8q0Z1EcSVwVUxaFUM
774QKuKf1zqdee3NcBRgNwpmANr6DCVaeyQMYNEu538ohGCII8vdObtUF7kBd2+Mr6rXrF36aKfy
l7sfD3j1hZdpodmqqSJdM4vdv7onabDIH5HKZD+xer6gJ0qfKGs3bpxAexgYGOCqB+nQ5yhi66j9
6gw/+gr4Nqgg7+wlwwMyNzY+6ThIDpAx6gwpMFL3plwjCCYByKUwr/dsoSKkeR5IBRmtGRz1t22J
gihGJ1T3alS8XevreqAL+f4OcMXN8SS0/w1I/uTFsXMDLrsFvfRVAmS/LHCANYD0SSSQ5Zq0F9SR
QK78NmcM2rvEG1NdAjxdx++uM4SY4ot3VOd8732haqQfR47dnzorULn7+ousgGufkfK725MUZ0H4
OII9t8CTzsirzKG8TzBF/3JJRitMwQh1wEpdGdnzhv2/io4ICAygT/YRlkRzeHAiwoo+XlquwS6E
gAGK0mrxEYWcR7pZL8TEM1ouR5PVrTG47HNY1vgK2CzdcVgDG1tVI0AtqSHI5htCZQf7+2iIQivg
ZpmNPkaf3DeG2oYg1l/mDWE8ebmNSHXoPy778DvZAVXXJwpzK+XHJ3GlrOU9N9ICxgyUvtbYIHPy
8dboJGtioBQg0qRuPthEKQ9ePyr4R085sg5O39IyXmxJAH+To2KbpvtPZY0hX9vzlTr2daYvR6Pa
xui2kecE
`pragma protect end_protected
