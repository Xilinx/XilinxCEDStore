`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AAXM30jx4LaZ/wmQSGZ52sWMTFCmaD90sZigacLWE1hKI8eSB+fwuyqaOyrCAV7hAcX5VNAzxBB/
WVxoZQNSvzj5S6MYBc1xBU3q3OzCOWuBKj5Fey+6U59/qaPMW11OZ4UVlJbzNCnirNWH5TGbtcRx
tLL7jeBUOKUW+UXQdx7/CqZgSDVbNs5NvYFoOTZERN8DOGYEB3qrdl7aPmgHooEDJnlwTY2TlvEy
1pSY8HDXjbGTWFfoI2MEl7+881YzmgRI2GQrZzy+J5El2K29GdgQAp7xNeqcFAgAL/kz5HlqobHd
2BhGdEtU7Nabdfi8hbr9cm0y1QIfT8pK+4bZCQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
ozn9cbBtCGg+bQGB+tl9qa+EWTWsJjqKP/uJZtHFUHuPUSy/s4Sp7WE26uu/pzFPUFZaM87pD6zt
287E12LsWOu0yk0RMS2I5G12PmfVcaK0RHWZa2ZFm18ShspORb6qQO30f62Oc5uu8LsYiYa/8xJa
ZLowuRPMOS35ZFHsDtsGm584UdrODdhc96qnfWXlsWh4gzdVS6tjy1BN8lnwkGA7d1ynsHj7hdVO
UaCsSTtP2n0yYwcKcs0He9skIXkY262nk5jzG0dvgWH878AHYuV3OFbaX5Z79jKa7Ib7crL2IPEk
YJdIk2JzXKlx8mDL9F9hotMOzN/oFkWxH/cF4vvDhRMFp9CvOvV27cMVt8YGAkag8aCKXSvJsmNS
T1S4gRhUbERaZuXnB6YtNVc4hwpN5kJSfEjaKBtyUGZAPngp0YzTa+HDFD3lG9HRwDpHX1pyk4Iu
UZ0+w9fi0jrkTLTf5MPmOJL8lnc9gWYr6bIeiS0+5CWmXV/Gk88Ij2N7toi3ZphbzeXWYDwt/+jn
1D3z54c4as8gxRlzPrCODNx68pQNXzpYA9URGQaoTZ71HttiahDdLT2ZOSbIiPyDPWKAyQ4zFhMG
Ijlal5mNrAtDJ3Zfz/iSIBvau/J8Jb863TcqSIfe0nh5O2mZfWvDzWxqKvo90SGMZYKSH9U6/wI1
Z7pl3QsqieU7C5tW1AmBj2PfkckrUQUgvHheiT6UZpkgBBlOGGuOwBSiErNJ2RB5kAjcxLg5fxdH
TupycuwXjdaEiIu+rZjcS/Eh7I8tTIeWf1tKfaMZPaAgbrDUBewvMTl/+RZuaiiEawZKbNGErDeL
8qWg94DvOShhrkhoWqkBlSUaQH7ThWP1R8jPGxxwBS75BaC8lemLQ/YzVtvcMAC+18IIV9sbdCAk
zOjG6JeYYSEghWjeQ5qeWdDUnIp2VDj6xxz5lbHvqe1saBptxff/IbbyoNuRne56MXjeL2PFyNzb
DTafFHO2dtnN4B74UGwU4cnkgiKqgZ3rv6aVhkhRSSC2KrRmurqoB16oWhv52P91KqOmrxNuzGCw
CeFhyD4TU2l4fX/JCm9C0AqN9BALMByM31cMLr8FZ30xwMcgmYG4OzCYBdaNyE4SjleOMeK7GyUY
cVOYnpDd9P6Kh05eUca77ZY77Ttk8xBIKhR6zny9PNVO0Mt1IdoFWkrH5KJhTRS2qVHPctQ+v3LL
QFJTDEB/u4cRgwdiV7uBXdKl2oVgd5UhajJo/RW4e1ez47ueP3z1VN0vfXL7K1cPJlqrH4W7CR4l
7Z/qTGl4d/h+D9JUDZZFcinhR1aP197y540Lnv/2SKYWDjOedolXnnCJ0hcOhcmSG6RNaS0rU8fK
45FW2JEgRxQKocnzW0X9uzLYvUDko6kN6GmFFfTqIKrdWAso3f3UQpn+fWgF8Mz2/8uIF4cUFQb0
66JoXquHAzeBgA4CLX+Kz89BwqNjDdFecESyDur5EKl07YPdSzg5rDca9FwubBMTkyX5cgvg0jhl
MI3pq8fzl3FKu+uVC2WOWmv3Q0tPO4+OF+T5mpbjEPReNeyZXPMZz2EVDMgmd8LBJWFuSIUZcgx9
qZZ4ooTB+LjEpb367irMKlfnNoSrc4jWdG4lopBooz8uME/4fLEkhw9yZRKDTB+0ZG5Ecij4S1sC
Tp2CFEBd8Y3SgWb3m/M9VRT0rhcRbg2/W5iM238RNjPlK0AFVYPzB5xowT3K7hNFHmZltli3rOb3
A2HtQ9zShd/i4/wGS/5r8wD/8Zk5IHN89wihGL3LNz3zRFTVGR1TvNP2fY7bwUwHBsMs1nAI7H1E
fdCUdW56PdnUfM+TTknf5p5/yo0nSJi9sZerggideXSUZJ2rcvn4PApWPLcRDDaCIajygIy3Jiga
P/TwvkoPp8V67o+utRjjhXp7EzPs5rtSQ9d5Plodz40RY5ioVPmAipvNpXXboglA00ZotLMOGAhB
nQ7WOnFM1WjMb7wlfbF/2CTwxNn1HBZulAIbOXQDyQK05C0DWwFNI2HOPCfyJKBRvM9jmvRUFTPz
we6LdqZmLw5FDxJtQ/xTHP/FYWMbZupGb17vfoeZG2i7sE+Vdso7U7KG2byxifw6MwVoFyza1fDh
C8zNKEHVYED2r5xDz3L/sGsmx11SIc9xm8rYWr/J1o10edQLMaUZCdZur93tjOxb30/vLa/JI2qa
cTBfcDAo8BKk3UXOozQ0HtXpHrYSZgSpcxzb7szY/963aHWRBQrQ+IeH0cCBD0YJWq8aClZXQQ7a
lZ0u/awT7X2IWArw4BwTAh6XcSRx25dbOHaOURsy5qOmMtHhJYbnl7TJEsZUBsEGNkeuabKG0sS8
PyPPvUbpmNanu79m8SoAQudf/bCwtFaQRqesLZrr9DH8xO7m8jjOKRolB5v4m/YlW5t3AsTAdRzs
OlIqdpY80Oag7suBaNks73Iuo3iZBdHkORCM6bi9Sb0BdUMAVsJDBveD0zMLuBO6ib2sT5WG90Xb
yDNO5kkupuuGgFfILd2KGy8juwpmBeaG/lSGp+Za4jZEjIEvvyEAIPHLnG2xLsHDRvsPrdHSV21E
/p0KWmn96kWgHYNAJUaChIRk/UIDLm1Dg1puRMk2MzzSIBRMDXiOyM2g4krP7dt6uThmNeFBvZR1
lGVxLRP5tabZhmdZtEYfyQVUcYx2HRI1Dp8nCXGbily9VEn0UxBk+bPqAOjt+xh/xnO6btJ2xxe+
oCPC/a/c/n/MI6MUtmVKbhxEkZbCPPYaPA+zZ7ZnOArOzlYyIwlBCv0IybwlW9qBobstMl6nCRHj
paVSjsU8laRkhlT/3hKyC++7faH+CWAaThxeADdzoClWJWhqPGSoUEx8gWgXj7CG03FjY/z9hO4J
9MxH7ndQbd1WvW6ZBrL565W0Z/neHt6DRkriu/bfd8PdpGEIwCLNNE7OkiP5acXVH2qd/y9y1tpC
BQxbop9t1ihuWgla00XdIzzaz68QPluGNQ2nDtBWdl/h/GkDeS2kp7mfj39xNGRNgSDKceqcC7xE
vLM0Ey9yxDBws2tl1UHYZG7vhuBKi5idhjRsz63B9+vJTRS1TEYj79d5LQ5jQZRFzqLGVRWydja4
q5NWAmLUYixQVb9Hze6qf2+kvC7OHt8s/B7b6VnA++14B8FDDwEbrF20tOr2o++cwlvws9rJ8tWY
7Mt8z0kAjIY0DrUGarKnGvIddL/VYlmMaFHtMUNJmMZT2FmU4pE+DHU1h8zjvZA4Lc61afMl7uEz
dGX+cd3BWF1xCqIiiWSp6fjMWOGAPsW1dETQ+pt6TU8lZxXu1lE3+GhD+Q10W6ueXjOmU1UEKX/L
Kq6UO8oi9bVxhSQuQZuLWmIfU8WGD9RVzo3qNjfPrwhA+oOIuNsGLK97T/KXpKYRvC0l5pZOttfw
4dlssK/HjOopABlaj7jHtSU2RdFtHkF22v32lFHxCUh5HkU4Tyi93VgC7X8YCqFc9x2QySvMK6hi
bBsjP6HYQkb15FPiG3Ay0ZsFdyrKZZMo81V4rQrv0hDs22MX4jyGuz4zRhpcX57b1Om6KORRr4Xs
EJdzK9JjHOwV4JW7n0FQPOpT4lrpZDbEXFUEcofPKi36elg1zmyPrIb1UgrcRLsSqojpZa5yMqf/
VmwmHo83cmbfL9D8byQWI3yUZUqmZtcqLyX/3SRLsrycmdqBkeunJxbmk9kJm0tiwg09wSuLiVZx
0WriPNHfs+cg5Z15vjL/uc8OnEMWV9+Fs54q0q6+GFbjj3P9MoJZTZVunlfCAVtYV+px53tPY42D
Y0Pht6V4EMUdUTlNOhh+9Rgo6711xHsJXHG3s+jCHXUzqK6VJU1fhqMyP3eAG4dY11IAc5JaUi8k
65mkHKyJq8kWBdLU9PgQhSK/oqw3m8rDi6rCF8dtQ+jkMqCglEZbbr4M9MJRFvyAWN1eZNWx6cLQ
7O9/+UaGriu3FfzYEtECtgfC6rstNkEcCB+m9c7rRrxreQCSRbsMFMwR3BDk/LRL//gXRvaBeV5w
7/a7MnyxuhWQGYTN734MKwVW4tlRLiaDCT/1KWkaKtdHyl2pb3gvr0f+TrYj3sZ/mideWifX/Ujg
ualtFsykNosn4X92dkLGowYmuAT15QELNizwcqiPgj/AN/CZ0pkebVSMkdeJVc2/mOO1juS8fBWM
hFxc1+E3Mrnv9kc+H1LsGaW1QF9Lv341GbZerawLWEaOd2ovXznIJwBJE2sJR7nL+3KVo524gQsV
zV7KFmfM9dT9/WhyYbC6lhGIHUrjFg/wflCzQjgh0Zuke3NA/ANuSuvzHg+NEit86wa6Oe9s3Tiu
IDhxHzGQLL1vu6JF448E3nDzJC9XMJn3EjUH9g9LA4GDPKyPFdDn/c+F4m9KjiLWcxuhSqOvunuI
QmOcSGN7m6cP9Ho0Wbas8sPaY6CMyaaJS2JNjdQ2qD0XZY6EIIrmdAlK1mldA0DR+UVtVQGnJ/JM
dwc9xhspvrX7NIPq2qNmCKZfHSst1CiVNNvE3w5b8DBSZQ/D1d1l235mGVKEDLcfoV59lfPfiR2Y
YD0dnavWcUumUzQpeGPDUAHLyqd1jyH08og4bEcnIwJo78AzDM9H6TG99v/dZ/m09sRdD36zO8cE
J3oIBxn8VPsm+oj8vQYKFltsyLdpW3kCfL+WjTa1etVnFkQoslWucL5hjWbR0cVm6cq1FTw7wzfD
lc+AlXJ03YT/vSH4mEbqr+1RIFoamN1OJ1uVnZvLU/WOv1IYYjM09+pnNEwq2DYzbanle8j+mRrF
8U1AB9dIIjmTLUb/wQ1tCRb9Iakh3kWxNxMK6qBkjkqc1xAjQZOXksKHkw4PwOmlm2b2c0t/vAjv
pTqn6BDn3eXy+WD2iQPaJgJT21nSfDainzCUrDTOXHMNW2BH7uGrYn4GfwtEcSR7M3KoMFQpF5SP
3og9bEtj5H8EqnbL5VOE+guQbRLPpLeyXNr6JwrVsMjuT5sbzZ1wN1GeqiUrz3oTtSZILHt5Kq6F
a+Dz9e8621Elmd9AZCiitwNEPIHI410jmHfhwHwn48e0qQypy7gYV10zGj6JNsJu4AnPD5rD+Maj
uJs16TZw76o8Yzz5dKxgQDFEZKnFWEzPkmPe3O7rX3zYP3iyJwbeiFMpnColfKZ1XvTwaGWKeAbo
+cUvhUmV38zWj3B/HDlytwTwXRJfuUdQqra1HAJ8jQAyfZadPMtevy7ICJoq3oUHxraJZmK6hZvd
p6qR5dOcNwXvk2o7WsEPfvPjnQ3QcRrI+3uM3BrALadJuLEKoeZd0eRxweioRzwmpkSPc0nzqhk1
2NQt0LwAtKkUkZq+z7h8DSWLsCwlVB7QcFInkc1/mvAlywNsiIzd7Hgx6KyH/DRRNeBpfdurkJ3a
p671JEKBT0/HyaYgU2xuPMgfvXwO7vX+LT2nRaOfFlmOWw8s6J5FWTAu6i20zAgYO1eFlg6tsHmL
4gVuqqrSD01GH/19fOpIeDngI/QLVi2V9pwj8OTfKEGkLkFlr1GecHmnG287mLsq8G1PBS33JWLr
kf1J7k6dfBF2C6XknFKTE1jns79NqMBFPoztagr18os5WTQBSDupmQ2X+KYEyAltylIoaTOEd5ZX
ZYzHcbni+oJJJFfQTmWsenzGRLshShM+2GCdgcD/ICNMeM/rla0picQ/C6t+iK7rCE2G+OqfdBBr
FFMbbh6sP8zFtBfq+Q+j8/CXOSsOgRYhVBWZKL7ig12dJYSgxaaArKwJi7skxBws3m5ZG9bM+JRj
MMu0HtuK/yHkkcROMeEO2KSMjQExlXEkJQpr+Rw+hx+pmUwZw51TZHlATXTX0OxfzfLsn6q84y6a
pUu7aqZqSbnqw+5fQneKijSHKi80I2nn9GQaWQhtCVANt+GDSwEHqmDD8b4SVeEOHMoQr9iLK3O7
3AYIjZeY8owPPluk+IxhxRw82IdZU9o69BFugPerPd17vjTlhO+36BQ9/INTkA09bmAAossMzzHV
UlDzGvkW83rhsLr4uaH7wh+MPptstY2tXuvFjxPISk6YnPlHCgD9SOKw3LLCzkSoLsTxIXmfx35i
SeV9ricAArhlaqdZI9qYl5e8fqCt8Gn3LMV86VuTDtWK1DcD0PqzixMkeDkey8dYEIaDbFUN9V+C
5u+Y5sxmd006QUpIyK8WHEMM8C+Q6pZrbX7McIqAw2wPrKfUhYPI5WvCrfPWTdZGnftMmafmP5ZP
BFHC+FD19rfFYELFBw9mO1zRQ5m6Sr0Ktsbd8LBd1s8nL6k3kxKUw11gkf3zb1M/4fYd+NkBPi4w
VJWsaxKDSixoPYbKSKCQc7NoKEd9OMHJPbmLnM6JyH5vbBu6/st59ey8XgV5WgwExW/Pn4g67k2Y
LkAwMxA3d9kqVP0JtoTbqZ3m1ZWiq1Kww/e78q4L1+24j0N2eLsYHNzuQyEofRVsNpksOGQquvIQ
aaMLFVBxemGrWjGfnPDeHkCxJ+XrD0LvTBNV3uRJWtX75YEoWD+cSsDqfna1vK8MIDuzjhsvG7ve
OsWzjoYoswdwZOZPPuDONZ1pjYYLmycnwkDiyDn4NHnKOIasdq5hGf7b+pvWmO/otik65EbeCV2h
lks5IP53NghA8pQRehJSp5IF4XUdXkxXNs6vrSRP6ukCE3suCqnKwp63FCg9U+U715ezBQlNUTT7
S0FEA1ILULtKuHKRsOyb3bGalvwixqPWuS4huB7g3/uQf9pBoc711vwV4lC3YK/v4f8zL+OqtB2m
MY48KwjgkXyIOHkEX+0WOexOjWMg+TBzX9JziQ2Hkgw7G7okqmFYSUzBVb9hEmc5mu0mhOW6qRqi
8ySAX8TjOIn4IC1yK4+SNHhi4ORK4qZrgjhG0QRS2WAjceVKAclyOyfAEhXFKpIr+DMBijEZqZcL
siWFA1RVHibJ+RpK7apz7dCHk2ltKRf+WOrZAmFgKUQfKVpPZkBIdnq//I3IQLx/n2F09b+d59/O
jJYLmHlWBbjIYazYuyQK3yO9T0w3VU8JJo5koxkGB8C+50lfML3p9uuHMZz+kFpoqGesRGWkiVM4
lMz4vCxL0ntYfyAdLZGW+ofyL9ZrTNhi1uNRHnB3owAjemh7r0BEWHn89962/kR664clRP8E7nr0
def/pFb728c/FyxjqnIG8Zgc3EtDQpa/OBARFRQcoiDVVj/Wxb/YTjyeYhxUmJ/8A6HqkfM1E8/H
bN4pOqCEB+jPwLsRB7s/O/2OuWMhgvmCKjCWkBKoNu7N98dUCNEOSgptzOoDdB5waPjAEty15D1T
5hA1DXf48wPdJJCN2mPMjgB94wSCrd44+Le7tboCsgy+nF5WC5uWcQyO3Au/QUeyhc64EBP74Ikq
v6/XXZYH8WnJRLGY/7QusA0U2EerQRA5Ev7fPqj0Bku0cK7Bz0xkmb1TL8tWne0lgrKWEdnqlAbZ
ebhRPg44kmfsebNWr/ujXVUqOBYuj8qUMXKj0nNgQn5jeE2XBHgwIZ16Fiju/SweszMm3g/Y1Tyd
wPJzZbwdGwu0x57HKlqL3WUnfOTP/mVjEv3zp/uXyiKyY4kLq9xkgyr8PO+hvOiarIDxGo/piX5B
gAJKt19Z9pXALx/6AhRgrNXV6nDvD1I+i6RLRnufg9j8x9aQQNHZ30RUSwWMKYi7Nv7/T5XiNBGu
U8kxD+fh68e0bJzNVUBPoEk3YP2+a+/q8L6BK/0JBcXp60pwgbll/Ui9AvmFq713RTnWI1Lo8fZe
abTVU+iKqezRrcjZ/VlaoQDX6RXKnh5RYUtWkOtj6OQcO3HrVz5tChsxezpCkvzquUj1iRh9N4Or
o+3f/INWMRB/PU7l01qra7UJ6On28/yJWsKnZzssINEe0NXxIENg7TTxrWe/aVIj9HvNHWBOmeFj
Z0FgLEVMJmD9sAJdbHPpy+CU2c/r28PdHvRrwsUwliJTLNkvHSz84+qGjzPLoM2ZDOQPWDT7NNYt
ylOy3HWSXuvCUK+x6/e1qKK/OWbqF1b2XRqdLZsmIXgfQhH3HElzJdorZMSbFTadYtZN6PBasPRO
1Edzk/FkHHt+YpDdfiKj1paOQnc8r36sUP8rXSpjxU0seUHOEqtaHyFbHRjCMlXUuJAFrJMmEE4I
J54QpHb+JjLlyHDDzAgEzl4NI+4sWbD8mw4HwPbFtpTNfPmjbNblob6a4BQTfubrcRRcIuC3ftfd
9NNMYjXdJVdG1DGMiQUFol9FY81/mo6W0Nxu+8sRT1hrjuukQk1HEFzfVHgy3i9uD5cQ18W5ck/a
q1AXQgOcpnOAf40qNjbJI90TXCfa2eJnwMBxc5rP8kiBdx5FTeWl2nY3mJ8IYVA6xL6PG64FBxwY
TYBYzUFI0Ma21YfxjA+BqnY+05Nbt+/UvtsACOkUNm61Nv+jM/5w5JVohZ3JKretPEuVyQsj89ME
SO+KkdCkRCBuGpxprNr+nY/eaUjmlx2wk6PfMhv7/RVJxhxqvxJyOYUmillWkkpm2O1pSiJGDTCv
sGfbIZLTVwBSpF3elLJa2kir6EmvgmWbM1dXPNRLYxBsKo7ttoxuln3J2G2tQFfB94e1Ul1ZCj8e
hInqHP0TjL0u4NzhrBlLAuzm+qyrCEgp+Pg91KcnBCfRc9IKmIzoei3M04hhLKlMs0g/8H6Yz0Da
CNoPeI1YKiWCdz//MW97k8rrjH+/JgNhz0orgwWwVXN6CAEh5K6its99YcHlaYXYO4I9ZnqYa1kd
v1OoTNItxQmD1M5kl6oCmKg5+6ovN0YqqGCoe5cAJt5hM6ZD570cuQpoQu+M4ByHyKixZtIsAOdB
PGjdKto20u0/fl7Te7jj9ujKXsOoD3Vyus/NOydfvUC7aPdlEZVyUVSzxXhwwljTNkL8xUvGz7vb
6pvDOWsuh4mSmzSsBhkbVcyljvpsFP7NuGMeR1ldZ36Ya/otw2Dj6qpJwvasOX86lpfoQ/+CFgv+
ZN5eU5N9BjlEZKgOWnZRg2k5xtblOpmwZZT4NI/4VyvOOjnMunQqszIo3wta/i/rffMPwWv2HWb3
QoYxFh/RS5Ogg8bvRo+UhrL/tFprRsdHOOfSZ5yu8Iu0zhodoYtUvUxVvJ2n1RkngTRxe4Hqboi+
35NRXFD7ih6QJxpIPSBhPvIItTs6eDEykytzJuhRHVILh+uvqDed8RMXI5op9/41kdmxn9Cn+Ewu
oxl6K0n0LzQ5EJTI9aYA5uhQrPyNa+bSOS1oqNdNMdkPZTwVgm3izwjU9WmvNazhTkD6r/M2y/QL
P6x1gEdHxnTqeC/xbPILFiC+GKbk00psPEO0G+UHOJvzUlYTZiZ0E56MIc0N/wWyK8A1AHa/RnzT
HqRoxcsjMMqYtGnOL6wzBHRlsmho+hK2OCrqpG6zpAT5WSqz/DN1uOraFQMAM5QRQf5nfBZc3oic
szg7KfQz/unuXKrFUck4x++mB4mkvks91rd/2B4w7C8Bgw7OMVqvzYzzw3crghmA54zRYp8y03tR
bAidEcpTo8iXfFTUhWQsjyXonbw5HLT1PnXcOyJGpgDbxhIWvREuTSWKjCK3tOm6iW6X9UYTlYly
k5wcUyJO1Fd0AdO6HKyQ6RsY/OysxdK+yLJamZiNBhFAbqLENuNyFyd9bftczuu8H3oXQOsPlgaE
+YFqRbUR5FT55dNIhD773jyLULicLj9D7niQ6YZluluq4FQ2+BR8nmsiN8qyevzkd4cMPBco5oCH
lupFvY3Iw18fnrJnOG3c5SG55qLnylKbkAE2bVUUVB0VqzE3GsnN2RxFuplMLUoX8pqVmB8qh91t
/VD6nC4pP4LHuupveLAk5tqhn3kfYNpwGVKHtUu/tpLDa9MizQ5LFAqj+vfz/hOmSMxGM8B1vikB
+a9Mz0fZSX650GI3RW46Y86CI3QJBQywbDjI65ceCr6C8kVG8w8mzAez8J7kpA2i8s6quswKzeHI
QdV8cE5pwPm6UwWJhEn0mTKeY+W/xXG8aNQLs+EBHyLd8HYD8NuoLUrHuCFeWHJBaLII9JlyBonq
Wx/Bv3toUXXLttuYqYBgKbjlphqCNl5j5qMCHKqN6BciT7WYd61LdO6UbuthkqaLQ/VVHhcaQzAz
NStY1BcWr3aIQk0rnCh02EDkokyR4OEfSUgZN6BtdtzGPqG/F8ltI9fvJXuwolGi+T55Cq9GcouG
XAUFPWl6ylt59dix3DoJzoj9ei8gHtltsCr6eE5CJIg6bHbm46rD0TT1gXV290LxnGbmm0RHBPIV
RnU1QIgXpK2DgRTNOZNWrDnXV4r/g2cr4/P/D8Ph43JWqCsoVIEa63gtRIywDKW8MSjiZrjv2MFD
CD6jElNQXwHITsnbJitQ3eMcIL76tzGRUuI53c9OSx2LGfWI0YaEk7bIww26w+AZbjcyMMsbf5oF
w/BIfJJFkOirRJwfRsilpi3eHs/ff6j8RzQZok8ZU/yBbSB6dG734XYfpWY15hBu0yOQfQwNS1k7
8AVu0BlBLBclm3g/XO/gQi9SgekWKrAVfwLbQ/VIB2RMBahGukoKrnkQiGkWEKKjnuBI80NUOD2F
mZ6f61aEULzMcteml5LQ+ARtd0QLhGeT01QYoRsbdqXnd7LCKu2bQjhKVT2n0mNLTwtYxLLbXq1J
owIn/sXTZb1b7mi8bb/oeGFKYKJpt7sz+sJOrayEGlb6yv4XtcIMjoJdyZO1wU7C+JkaortFoGvi
Q+YW5N29V30rOIdzxR8W+oHDn9W07mptGqmq5MIs+ocRTdUNTSxgHxjp5KqLcXK5JqHvQC1PDOgT
3M7fWs9P8SeDvcktpYvtoolOE5nQPclVhyvHbUuSiT+C8tx5f86QUD7QsZfYMFLuhnsGpJ8QSgP7
0haD+D7fkRA8LNZNjEPXIWCG0BAiP71PX0uH+92pX6/ZHswVXVN2ZJ8SCwhCf+7WzDERvvu0Lw+7
dWJOsDBZgO13c+2MTdWrLEbG6S7IWiIK+PnQc3BLfif0H8WWPlJSrtmOpLbc4V24Y0a/+ZVtz59V
mwTDb9zcBTtB0Hrr79z6vclCXVA1WqcL2vxXsujyzEkoFsgrRDCiVsqkVA5jwyo7oyD32yLvbU7X
RqmK3VW+CBKTB4awek4b3KEQdrgT2WWb0m6tCZEwYM5GxEJ91P2CdG8b0bPKRlScIht6Np4jlyoZ
Bq0EaZGQDspntI/t4upGndhnKe4ozDFjSqjJdBjvAgaH0tZX14dT4p8yCmwFxBBaybxUB9PFyGUg
SRU+o42WgbNIW4B4cAjtnmpCZAnrhWL0goPh23O1Hyt9H20vhDCc3OPGSMIBncf821cBzm9zTHc8
yWU6Fbbz7eqyeaM3rS7G3is7yiEc4pNY4l7vh29t0EWutdyS9GvXbNprfKjR9PQ7dLic6VbTPB4l
OBvH4t+rnOMvEkpV7jZpdY0j/T+p3kM54+jgjy8g2uzc1yZXdvSgUkxUvI7IbJ9SmpWgnF0P4UB0
5znmkHTtjOkK1nu8PUoS+vO1EvRMueo+GN5HNj1Ie21jmEM7RvqoMRkr0pcvq6y+eO3QAp/HzRDY
VAy2sOKM7YWEo/MMtd8tUqDXuOryKAfC7eX5ozSdg+axuFpynDAHjgRJUuIZDHkJicgheWqyYDlG
/Yt7GE2mq7IZG48wPY0uDRT9CWZixM6QjXkvXbEpA24PjklpRLz8DNj63LHLq3wR6K9zkY1PSx+P
Dfl+H1X5VUKm1VYtMGLeuQTkIXjCGSAILagqxhCV6yoXNxvDrh6l5/NFu0byQ0CTrTrcggIjZ6HY
PLmaiEOTjyGpWLZcbO63yLi+R7LL2H/xIX2Fum6DPUBlu9BsTOiqFebEZzkcSMH/EjETw2QjfGO0
u2aCrkkfdhdO5gB+tF+feLM2iq8gfzF2hNgdA62eUfNTS95itRQNNnlT3eYUDuBrtKkRRcGsbP4p
Vf6VWz9oF9hpLdCJ7dEgg6dT4+W5efAmtkbbZKlSUcfcLxJsA5hBiel+sSYT0x0i+RPfROIgFC7v
IHDz8LietzavU9UgXKAgBgrYJz3muhwd2oQShceFpNVcf2BJ8J8y1BQmkju+2bYrLXHIuNWOIww9
Fr6PvqKnPOxK64vgNIc5+umX4rals81BcV+38ghdNj7tC9gfaNv7Taeg2D06BAvdJyWBHWu61NYg
qBNMLjsnTbg+7q4WAv3q72OvSfLeE8u94rz2TJwMTlL5LkFGDA3PMWDlG7t/TBuUH3KlMaSVtiNm
NFprMHR1AI0HqvamqjmzZ+uhj+VmsBPzp+gC5D/vIeGr1RRztpaesWZgHNNKHoyrg6bf5pZMb5gT
Cs4Kyi2UZKI0xnnF4fpmk++WFfofEiItRwlf3yiQ8FUELm41lXKdPb2q/OibbznRVq3t6T8u3J3U
5JQjuNck+CnQZz/STLih0dIOZl5R56fxUyVV/lLDzAeA7NlhGbuthMZwbMrpbGCkTfIdbJd8viWg
Qcoxuha8Vkeyl8qWZeeHV+jxxmOyoT8fkkEQgc85cB2OxfyIR4+NgnGHlJ04oPAx1zJaVBYjTaGw
JiQuzVJ26tksjQ/lK/7sPbUWtc12gitqO+A6nPGSXLUIzK1NN4w4TdIeZ424olOGXgg5HhFOyWYP
ete5aIyMvQDvz8G0LcR3ZJL5K1HxmOGd2gc3eODVNGLGsW20RHv17gJXbKNu37t8ETgoLx2cFX6r
6Tr6MjW1v9jfhclgxVq6hHjZr89faGCZkmm1RAoXqA4+Uyxr1Duln0mYaf9nuV4va/4ZhnHiEQkg
8d/78E/ZGCArfTjM6ITT4WQChkxQa9rPvXDjZ+vuX7QGWkAs2uCHkk1KwQhY0+mia31S5/fVVoSm
vZ02jDncpq4rdKsZ89MZ4kR6u4QrWy9FZ2rpQ5QC2axMyet/iOGE3AtsdhL5hOkmC2QSRz7LFg81
81knOq8o+8N9pkZZT5Jdyk6oYOEYkSDdDODEyfwzmW3Nke+pr67r/kXBgANpS9OWdAraRu0PWylw
19nzrBWuW+UfvZ6rgaiD+RxXnGlkxh5o6/RFMdh6Nsf2ZuOFnixvH2623dkM4Ro3Jv7k7jE0G+hC
4cjmAux+qHtlC9B3RY/Mfw76gZYtMkmbdSvUdJxSicbErI2dkP/vApoVsPrzhyiy+uKYVZjp8Uj/
qYBvPFXSIJ7JP+SkuR+v9Wua4/ZuoyOTOjPnKLTXFgeP7m3EjkTkrx1J07DHcL3gU1LwXRQ+6Wz/
Lj2oshx9WPEZ1mPfom01hL6R1w1/fOZp+GB36kejiaLsJS5WVXQcN56wxbL0S7FKr6ediJzsjQTT
brFUyg1Oy1ZAA+yPGgT3hffuSA/l/szZaIiifai7KeIc3Is/5Ir6h0NnmlDbpHgAJ1bn1J110u12
AUVH6+RBZ2rKVY1Kpa2mw+uvRkIcJpJqrPPFqerZvfZN6IXkuiEFn6fdq/OPY5jge0idJGekmJ8Q
uXDpqW9z9ToccBiqt6W8Ne09TT/wX6+5hYo+9c4I1+okCQu8mQ93UGyXjFfN8kw0p0gTQE1Bz+Gk
3MVLygQdmo5GSlFHTgasV5QAuzIKoiVPQy2zmbk7silZKB3bDt9H3Xiq6hTHk8eNEma3QvxyBe2P
MdMZDfheKF5f7ORF2DfbXFawNNq3xCImHEwEz/Wu6a/tl6JKZgpmmOrBCDKvZmbVTouLd79ndsnc
+iHIjLoiKcpLD9OLOKJRvIJON8+Cj3hLk5Agxw1zD//yJTb/2oTiQEFXBP2nnzcYl3gCS5/apNrz
qK6jXNU6203jbhy0bLbl0Sz0t6f4Ml+TTzLznoDu2WLmHdVrxsZN7/b4nEgKHh1idzOQ/QW8IR9u
2eMUJOT0ehXOWOYwirD19Oy195UeVd/PvF9uhc+mphg7txzjtXljbrYspIJtNLH8pTKmT2dyc/bg
mzRuEHoSwYE6odBu8YoWP1rLmACN4Uo3fxe5CHEZmZYXFoqoijivekgQhRTcv/Kje5AopNxerxad
zGgChsjGbLmJoJIkAka2JV0HzW0vKUOVMdkM2+8+d/97dN4GFnbW2tb/8whsztdXeYYLKPAXghGZ
s/hH9unibSGGSwa/QoS26BtDhGJs0SKA9RStyrr5ZayEhR3LlCmO+pYGMCCDjn7FvJGZ8l63SwyZ
Igd1/Vg8jSQpB55gzi428uOjv2NZsCAwJloxxLXsgmlCRLUqS/onUCB15FCG8HbNAYUIAj6EAGrd
+L5me5dvGYN5tt9uW4h7vMWoUrL41TO+D1SlT6VIS7zBGYTJTWwF/jvOlVKVpH1DuDepNJxeHn9W
48p3vxWscs6FxxnMvRY/ito+3wsuoatZG/LJtkBZYRAlDesVUWn5t9/Q5VL/AbVDqINt7vRHdrLN
wN/Cexj1YKCBKiEkGXCCRjf9LGwJlTRzmBLuMxoETaljuluhWs3fssSclhADAs6xoP4mLidkQXIZ
TrZcaYh+O4yY29CkNpt5TSzltHOCC0Vh8s5syyfFWuL+vpG1egt35YUqqGltF79/e5BuctJQJu02
76KXEs1CyVdBG1hVO8r+BEtF8LXx992iLCnlsHa6SbOF3TQqiEhAv9WkrpAxDUPFJy/Ov4pfNboQ
a2TFaTvUn+G7sNxc6ZbRSAWRXD5Vl63a2dir/KY5jmrmdc2sYXPJF07m8r3j08CAQrsgAKkDlWCB
siR2wHSVglAyrIdW2ZVhP3b+H4roiC5Zy0Hn7iVgIaFMLFN72InIBTzywT8qFxbDl/wn9frl7sfc
U4l+fDEwONBbmSvJAo/vq5iZZB0+oEsUlxFrRf8YdpJyF9ors42wP850+7ns9WQXuinuf1RDmsFc
Ntlh63fpRc7xbWpe9SIJty09D4OwzyANapd5RFrK5zIrZghtcFoRJI6kw+vquOUcOZIovMoRIyTF
AJcT0pKYKesyAvGANp6W5xlKPSEGe1piW1CQu1mRHH3wOiWL09bX8gKRDYQ6YBP9pd9dAy1VnchF
xPpal8cy39KAhZcN2dq4/Vai9Hzk/L5Wd69+A8fx7sAtBmiqnnTVc8E2xol+w4knBsWBP2Jjnfye
AkP9PQAkvVEzAzw1O2XU8WJqeHrLcn1k7ZeicrFw5yzeQDDMDYagUEh1T2eDQS3Bpo8aa9+eJlDS
zDA9JlWXi5dqZ9vonfDj+yav5afzBYLUmiicX4A8ngboWz1N3rR2KRXVm0qRw4ovGk3Xoo1YXeel
XBPAc36gg4tsdeUBr7V2UT0qFRLO7rsF/g+XrC056Kcf0+Y3jQ+A2HZDD5UqQF0ldkFCmnenePzU
KtM90GpXa5iREnrekE+ZOaTrzYCQ5ygLhNsRlRAxxxMnOPjYe393h4o94ztzpSHBKCBNVbJskvtP
HJeDJGvNSI74U3vn0NQPDrGTse4R3ugunj7pCZoLJKHyPtTWjNTmbMgfs05mlvK32nrra2+J9DUX
q5zPF2kdj54G0cLmThrNev8YQJa5KX0YdUrfkaQr9UsUA5qRSIsNSlbDt7r1r4xIAL2vImmKV80L
pvWPfAOdQ0B2ZwHR/+8JQiYL1O7YGO82kMtifXrCA6M1QVxohB7gnJQBeflT/xn0vt6AYydlff9n
8DnGuNe3ZaiUy9TGB5IauNdWrMQsOB6QlET6FYxbeuW9ZGSmpEnE9pPlt8fdq/Eh2IGTTdhxSNxa
w7OCnyCTmW10Om3oLNku7qgOvluCUGs/LSK7zCpCSod86Ys3YoMEIHTwmZDKbEKGPE/cfqiotjBM
dgc0++iRxznm5n+C/F558Ae14m0208mHNsrpXjQmy6AnJpWchDxbdJF12ZwYlRCgwxHBNolmytmv
mY0T2D5Vb/3R54vN9Ny33JdrRxkx1bjX+SZXcEvUe4fulrMQukRU2UkHx6bIJ/9sWUSjopGhb1KE
jHx2qM7ceZhOSFdDuHfywAnS6qEC4LuXXC7C+MvQt114r8RqZGDH4qEiVQG7+0fpPrWER9InKUc+
+BjFff01yzsIHZkJLo/+ZM7e+5RUSeBDHbtavvCmZpPHtLBlYWROZ3rvzRwuu1e/1HE1PpFL0z2B
fDUg8mtmJLHDZzkTtN07wM9cwIHFJK5NFoWlKpEL4Qnt7zYl6qAHa5HDu6u5537sTaFZXqrpfGkt
yF1F0JYjKvcxaV6bBzHhWRTKT8/91/SFn7PEliNOqQT0vJdmoDeCK0XztAqfPT9AeY+ksOmIZs3w
QY2buPRxdTN8XT7F4OB8IvN8RF/HFZ8mLKRIxLlUWiVnDWk8du7mG5OMA6E9NcpH7cR/eGud4hSQ
1l0ecQDaZBwf15Oty9MniRh/ZJ9csQldv2bTUBLegcfWzgQ+8fVUlF+iWfe5jqBjap9nmclmFTYX
RvFI4iNshrNQmIr1liR8eHOYy1C/Tk9H4cZApK4sTvcNlJezOz7kIlj8bkA+K+eWs5IIYUM9hcF5
orMZsHla4h1tTB/yw4xtE7R1yOvGrSNFBMupEfAPJIGpP4RCo0iVrBCjJBqMFzvDH1SnkQHRK1vu
QK7ECAbHTgm+0ulqo0ICUKUGtVl9PUOxpqRrCC+63QKL9zWzc1ccBuRhYABgamWExRZ/SL9GITCD
lB3iAnxwyg04jUyb2WDyf8hvrhIWjmqeCrOtqsdWulfAUOEtt/eDNBzI7lml4vidudDohnKteEGV
JAyUwWeGDGcYFUnCxOT6A1x8c/KdszHJq7ZofhY48rNsEMgCEa1Okw2Rn8SjJg808zvOfvxf19fQ
Zw8bdmESxn+/xqoFi9pBcP2e/E6T9dfNjR+fWrBc/dCDnJN/NFswzlE6K+JzjT9vr8VHOGAj80l6
zBXcsCPuHUlTweBxCsqKKWAVDaZgHDdHpnifCX/C1y0o7VwqyXxhLz0o33It1ebrBA7JLbhEKQf6
R6d+hqbkPmiHsjFUs/jlSoAALEMapZADb8cvD8fV9ggYD/NVFeG2eDxIuEnbDpXfP5DFMTjKgh1I
4O10BNlKGWgogozAnj6cBUx9bbrxlm12tNzqkizno58GiG2FykIqJ9p34a7g/vB+S3aKz4N/E1MU
dS8lgEO8iUWth8cXINTkcSZ+sTl4IaXfMqyClNBGB68CURQdcAHzZqCxELd//w9KKuVWOi50NFUe
wV1vVZTzMi7YPMMY9Uf646YQFa5DdJqa7mnBe1F1A4w41EXroa1rEnKRuwf7pfUAjsqh9NzYz1cM
j+l/l39fUuVU7vs9M/0dFCsg0dr/Wdss+ZYk1zwsjk06PxZq6CMCGCHEoAnRXHRFREFpBnjMA1aI
Ew1rNOlmbQqO1z5qdJJPmviZtXTIkqRqvXdHOw2Yau0pmJGB3oL2H4BCZraq48Kied6TNM3jAKuF
rTrKsnuChNYvHtDE1GJcvO+NFZ2R4L7Fw+7iH4TGlRnqPYwIAiWDY6C69LzBI+M1qKztra4RjCGu
alAkGtASxrINaDoDsXqVwZJ8nEVhEKOsta6BcM72ThXMrKk2IBfck7JZbYb2a8TrOxzuVx/zYPOB
GZdR0ycgRIGHJJAxED6gfLQa3lyMFEAWaaNlNbYXK+r2E1LUk+tWBg09a1wPEniQ/svwoP1HRAZ7
XcyMIDZdkoO9wOr4znDvFaS9vWZXyjKdAYIIIkUF9W31isVWBMpK87dnDL7NiOKCqY5kXnGUZGvL
evLtxwgRxa2OsWpaGx8VSzS1FeKFesGjv/taL311Yzv3DEr8YhmBCqUikwVUmyti43rKiMrkgoSu
x5ystOcIrctUxdg1DiPvj6jgN7BY59g0JRfge3Nt7mAhsO/9SboUadoU4oRqE6A7KH7hQwpdXIiT
FAXwSOeb8SZfXWC9BWlOiVcUQFHeKbyOzhI1f7n4kZ0RFApJJ4EJZUihtqYUY4u8GibVRScXksqi
igQbm2eGkvf4xy6oKuWVDDkN9/h7EPkcszT3IJ00SyIkEkibJnhtoaxd2EkJ06Idzvxt00C9z2U9
eWu09Kp1dZbrx6ycZYvDPLUV09QXVEXMkxVg3YDpvEPRV1vrsoN+KGcZRuxO+sl6eWHLsU/K8kcX
2WrkUBXA3jrxSA7muMRzd42VqbN0COan8zN3HWa5QEZRfYvbw5sZVk/4wgTVl3u2ZPvF++VLho4v
kUdT1p0skuZGo2hnBr0EEhtMnNBJ6cw7+9uyvh0TmcmWdJW7aOF+Dm28CrdZ4i3ST/L5sVn4UN3L
j/o+zp7+fwriuuzgOrg2tB7gjrtL2JQcchsdZElWAKTVbAr4tScQuKItWdDOEJptFgj4l/zqbJpC
oCxzKTbWp7ubwHKl6GZlRpMSVeYVZp8VJypZxZTImEZgx7JlnYD4/HJoHl/qWGw0o+YNL5fFh4FK
Tkhbe/QkMjvk66rMsPBY5piy4fKFNDv71paTRfmgdSiZ/1fC/hXoZGt95GgBDJmlUTri/EVSF3MQ
JRM+E2ndRoJXN0U2O7CqxEHf53pRKECZuIujJ4ER/c3sVP7hxNUiauUBobYnG0BAGs6awqkR0NUp
Iz5gl2bAjfXZ9JxxG/BjgYz+jvjhNj75FctEXSFCsY5llHR+i78/RhV7z2nq2IznKCUHU2EAmCtB
BSXv6UtFbbrb1ASM/048c8SLCc7WDpvjqy/vqUFJXLup6bF5DXWqhG1bBZyG0g77/8uQ7NISzIf4
Sfnfs/JgylTgeQsbFk82ioRgUJf4fU0JQrh4fv493NvOqvvac/HGUf8kZmbso3rbowuljagk8JTm
2c8LCmK3q+7aGIw/tiBU6VOdInaPzw7ukojpc2D/KiiLoIz/XtldcxrOrWw+k7O8d7ylLrMwms8v
v/kAYDNfVewmkRwCu3U5wSzNcO15qB7GvAo8EP0edkuocr2Xrq3Z+YyTJEaYnWr7NOvBgAKAb5rf
3UEFDSyr/UMUFJRpj7leoT6ZPpxX1DStGxf4ilNEoO43G7FO9OwQ5D9/DI8OaAFaCct/3n6imdEp
vCgSVAB/VsmwM+KtBs4ofhY0WCsXv8pE37GW7x8m3pxUqGzeYdfnH5RgTHV9jpALG63Lpfzqme/q
NY8880SIV17gFHW+RswoxfgKXp7T2E0KE1LACklT2YDMETS/lRVJqj2cGPL+0eayhenhXDZVH2Ac
ExtRY9J8gzj12m+LYCuSiMTJdfDHeu32McbykYA1CHWmN0jQGuPsJOvqCIf6MohNhQwsogwQ1c/7
aePNv1opZy4/m4TxYk3QCvIkLmgWk9wnI4bpF9GRNQSH124uwYklnsUbBotPTnd2Mj7G3XjwGkNe
ElMCvLrLDS2T6wRaIrnYS3lDkSsfVLMxUXAyoNeH5mJAVAdUDk7b+pNrzXIagbOuUmyIkOY9ATYa
8NzFRmc/supVVY1PAbQDQGpcgVksXb8QxMqrnK1tTJiiB7sOamaGNZ3QeBNux2VDpjtkrnTePJNB
b0ccvfhjd1TKU9pgUqacMk96TDOi1BJdYw2CcA8YHTkuceUUJtITbdnVRCmnXngLE984ZR2oVtrC
cQtsjxXRaSPpJyObX3A5kiUnwkU8nPr7qbYSrowJtoVsdQxz+TZ7Z7UUUmbnvBz4JrbugJuQk7hB
YVVfK+hSNNET2RdAL9zgA7XnrkYohIUqlUA34p0tLe8Va4bdNtqGQyS9HbpkhzuwGUy5KorgxgZb
jNPXKasoRO77Z03uknYeGnz//JqzRhjq1iXQT9ohmMwR1GdJXEVh174hxXBeWEAb8GtqYMFXv8H4
kiePgv8fzB8oAqNFh83GwzBuHMHkkq8goAc98GgpjXa9UungLKLRxWT2JxKo+Zuf3Lmk/FgXA+cj
aTHYm271Q47zwzgUdBHr4WrF2eDdLyC5Uc4awAB2v4ZAE/wUp5fa4rNBgeMVcd0ekeZ6kbnQPdtJ
6mMbhyBeKhatp4HIXK9iHbaS4FLgi9AwgD7+sBWAPkKBo3PCocSszIs0qQu2/5+YyQU5Ba5opH0w
GHfTTWpL8yVNqzfB/7CQMKEsy4xMRc1wGHhPL3pjGqoORnRDgXp2do/FvZN3q/1MNXyBoNTutdVL
CouTknSX22MEJCwwKELa8KwXnCuy8Fb+JqBMporwzkJ773JdzIy0BO7tlSm2upiPciosX1LWhSUa
0C5j8effi5l9nP4batEkxz7Fs48oflahVumGxYsXfJ3w7r258JVMHMr/ZewAL3ppOHSntNZ7wNsA
bMjRXVMejrN4roclD+pvcdZO6L8QsurICrSv+3IPsrRJbjMwR9tlsVO6dB56KFEZhaHhUDFW62ic
sq9slfHtCwIGQakTC21eSLogTj2sWtNojEDabgQ83nc0C99eigJz0PWokuorBG47oMEFNfm94BX7
iSKwYoe7l50Z6WcXZZJADGQOvTCdIyUH09uW4utLBAjeg49jXYGCCd2TOrof1BcmB91IDC9qW3ur
Ca5BjK1vso4y2ufU3EDt75YunqzRViNUPtA7D1dbJIzm7XfYz2Ri/ixXhzksdaw29X/qW/T93eaV
8GJhZIy+33rkU1pqJvC7a8m6xOQ6IjYNnac8iD6YIJU2azDnGO00f3ZbKtcEG9TAnv6U86TA+k9M
2d89vsTX3ebxfjsJXKegSORKTtcjnFQj3wWUBiegT1GLZUYE8wAeRM9gHo8W/YjSnDz525hNt/Sv
o+lzfhm0QxXlj4L/uebQcM9vJqMWgVILvebWPpu8M0LUuO67i9jFtVd6A3vsaAACbsf4R4ob57Ll
smquPzqWvfvlgqIOcHjrnRqOxzSe3ky/Q6KcuSaD2GSU6ZNk4YUHLjYxr9H33EWWHpABUmySln6M
l3K/XPfd159lPrsWGA/rxlwXPMS8jPsPiksG55XXkz6sW+4nz1+MaSsyIqhsU1ESdshA/COFP5bQ
aVeUrFKy/QMSo2YXCuToariOILcPmH1cr2WYRr335o7mLMWBAtWiSE9HeEch50Lq64agQtyT6dwh
Vzte797UEJG0JwnYRrA2dZeGJvJLC4dMNKr2+0ENF0JIqLNn9XYJZnh8HIhOgCPmp2hmlNV8XAFs
awtDwVFEmiWb3k+vow9hOB/SXPv0FS8yPvETYYle3WJEVUjhR99zVDQu901bJtApB9EyTYlMHDdd
+8HGh2jw7wYIQ3hEA5tV0lvfSo3BuOaazH2kMiFbjezE3F/SuDvcY2KGicf9TQoHxl68hLd4VrMx
tkfq0FZ0Kr53ciZoz5N0RkJzd5bvw82U+bExOgTea0Q7+0B37p6RNqqC83YqRW2X0UMpodYUso0F
YQQLyGbFNfLG07Acplh+uqvNqfee/tO/QzSMCx4fNqEo8IrYO1VaseaOGoK/COKPuReKYvj3LW3N
A2PQDD+5VD8DDXG+Qor94WCBt6fi3MKQbSrLvOIeq3/j1CNrQ+g3lON/WGr52LFPUmp5lSG/7X73
cGrCSEwbIMcbOPTst5qeTCRVdlY4dfDsjt9NbuDzdXBwp1Y4BxhmpmcAkvnpDVGmgWJLB9qnHkIl
ZBRGZhxk6G6CkIggqJRv5FYGdYFKKtvoGmDjfSO6Ih1a6lessPmsyPHjcj3mWzI04+oFd00ZFSpH
7bWlYW+whifnhoyteeaNKGd72RfjyfkOF6RVo6ElP4kE9jZAULgDjrhISixDHySk/nLnoYU+9XMa
ALlP1FNmKkEox5xsQGVEBP3X+stukZBHlkOaUfiFZbFLGDi/hznxfM9mQlda7SZQXs855G6gEiK2
IiiW83cCOhzOhfvB16z2AY+F/VFe0FslUmEBcmV75e0oCzdhwImLS/F7mBFM4PCShXTmxbeJlaj9
b4iPijJjBMuyD9jDp6DFTg9f/JBfeE+daxWiYgcOPxgvvyFRxCNLnYucOW+ZznXfle+OhsvZafsR
mcjv+wiu0cnTrI2gBXp1KIM8ilhluzbaG/MzIv05J+lBflzshkRDTsLn+g4dpU8GhTm8zvqonj3W
SK0GGvz1nknNc3qj/pnvGdtuQupmvu8A1XUpBd+o+jIgvN8uZi6r4ZKvmBbGvgBw1y0HpzHB4HmG
aKPV57v8VQ7GpEOEwwptFrbCxhHPARQa1GUojD2o5VAAQD4Ii3N0HaXAKLbOGQ98Wah097ya8bEH
NSLAn0SDOOAwRMi8yW1OztE3WJguIdbuFw80dkpz24a7ph+OwLmqWJjkJlFXpyX0mxOfu+LJk7+w
wDiPc7DOJLK5fsHTmoyf6fsGeTnsbzkQH4TzG4k2JWnqNSiVqloMerYTc4fLdoYPcDt+b3+fpMtU
LMOCbO2hwKCXAEqru1O+7IP87HMrP9w+4nm2wzTRejRId8qTF1RqHlkeA0FVRkhnxsfQaZB0juaL
96Q1Kk3gxFNPj2cA80P3LM3osTpGq1Vt2q2zZ4Zkw1+6D++v710uupQxLaWIIub2Go3oC7oZrcrj
1ZFafHkIviGnmAfqRqqzlFT0Rsypjnd8iQ6nuW3a/sTEHL/wgFTvdbV8VUx/nloze9w5tvbu50NG
CQ323QLyvrin89hdoP45C1X7HZxvjuGFW+ujfzAcU3hqj4tEBeR0buDSYhKn7C+aKV1kImAnKvC7
Ns/ayy51zEG1ZG6fQA2nIVaQcJhN5X9uSGNY0Tm5x9j8qSUD+qVgqd2L3uYRXgwFRFRIZio7ou5m
/lHVz3j8yuJoGLSsRQM6IPdb7HpMpfaQVtnZfcoHt+tOVbrJRmH2glMW9bvsI/hKKIxRL2u8Ohx6
7OkmKxxnzw292r34Llkuy7HCkp2IeXQsJlumVl5C7ai+Zd6B4HqZxaHokLsyjWetKsu1O7TN4vR1
zux9sBLkUPrPWHlNQn3jUHoeCgIVHGLc6erXgM95EZs8VeCW6Ve8dQuhKBcplxXMtGvDwLxnz1Vu
KUtuiujDpwH00kdoIFW7FPxo2jOXBvbFoByHKdZi9fp2C8FXMmwtWF0AkuvyILOgqkcreO/ZJtxG
RsqGsoFrjbP+B0UwvjbOHSy9580yQKdiUaah8Vz1iHmDLCcRE7wLHLdZEp5bRPsiv83ls4QkTJwO
qTed0O+I7Sqp56DHX/GNQh31p+B9q4xPCb1P6JKk/u1ivhlsVuhj96FHdSdpUipZbnVEzQc0PXH3
b0JHeI9sfR9KRBWgGQ14kszklrKfDXA9mn+2CGjzOfYjqbt3Iyga6wyjQSmnxsTnl6llGeDuuUaO
sONlOiDWlb18lAwCmvJ+X+uK0pYCl+VmgwQSadOyxXTeHeO5QRyOZ20+mwbO18DiNBrI7b1OSbXr
TKeUk8RxV4KR9FMw/1ICNhi5GtXYZjLwLnUcOHCdi94K3KFKo6BKCQXrTQJ4Hk3M27VfVRyEXdYn
b9MbHvDRmCAS70vPXmD3pF73xyP5+IOlgnCNFBB5jUL23ot9wXprgZ32ngPWMRWAaoD3VASAGDpP
K4kJpqoMoqpfBWEITaSWqRzV8N9+j9tMMkutw96hpvxW53fD2VbAw9rBuQTimpKgTaOiWV2IkyYU
u+PX4yvv79+nd/+89S1rkBhWakJ6zCfKbHw8p/1NF9gt9UsUUcQ/M9UcRBbQ/tw+BdZxE64DmQsB
8ofWB6n90vfdTzWTeUstfaBLd7HPU8ZbxRGd/d7YZ2L+ZqZuwDRLbye0iAr92Wu+q0NqjsOso/8Z
qEFHW8dqusPqryXYe5cBk8GYqkLBre/c0tdQO58sa1hSLc/e/JfsPjymJKKiW08wdbrl+C995+PQ
BQBeW8vlZP4oPY1gVrFvKVaLhvHUnskJyvtK6KsKdOgwYBt+fY4h866LFQGvvVolFBuFkqPPWSh/
EwWxr0kQuat/X5EeqmAa4yz97a5w9z7nG73i8a8u7fJLA1gq/5TQ5+6gjflego1rExjDj+IchH63
3/xMHK3Gi1Iog06ql7XxHrad0j+a/Luu+JNY0JVSn2rIXBhIuw32VxUssklcHh9v9soN+lBCTIWs
RZ0KOvluP84Q+sS9SZKUx9jgLHsz36n37+6FewFRTLC6pUDCiI4QpwU/nB7UbH7YPjheC9HuZEqQ
L/sh+T6qDCv6ylvzDOTl/ZzO/ziKSuBO6nUen2rk4aaGT3/DPseVJa0Lm87JX1/6apGOgixPL5gW
CJKU2WRT+ubZ6mjuUBbo48x/UCgi5TLeIRTgr3By4v3y/AxA1HxbeJ/oDnMer++wQApOE9cF/isc
y834Yqp2UlykSxjXgAnkyo/mlDrqN9ZaNm4Br+rMza2Ew99uC9zIHNzgjmj/kNGpNERN6dLN6lK9
Jlqk9zg1ixwiiCoQqjMoPxpVNTSOly5vFNF4pl9GrHs2ic/XULpP1C/TZs3QNwkXl97yxfQ+Gd5+
tpM6FfpX+yqU6KE5N29yF10x3bkGSKiXdXHITAcVPsDGb8L7jmCm0kRGjhS+F3me9fCymRV5MYge
X5aL4RDIvJnUDcBXgdlhEQgQ3zTx7hE91hmLO9w5oMgOutCqRKVTtqiMHGAsWvPPzNK0ZZnC7DZj
ubQzcpBrsJ8TUxB5r6+C+DpZ2YFrAckWXUOM42jGhtYEX+118bhGIgjGRa8qfsYwvYjHR7JnWLL3
5STiLCKvljdQxKMobtR/S5Iizjel7aFuuMS0yRpw7SXcUjZbsVoAxI+mzj3iML+xXJaiJMetGMHM
E6zrsjzxOKozfDdDMdFcDeOAM0xd5mmtuoxoDRWDieYKyyi0ZrxrZCAMUbGiVNlgjZbYO0+MbMMF
oGWzj1ypd3W3kPey646PyPhr7enFV+vuW9r17UtGDgo7s3OMV8Mngy4lylxGtuAkGvBSsSUWirXg
Nhtb3YzNvf7jRIR4guNsTTf6ShxDkHKYIqVQYaH3fiqAcCK8WzpdBCH0Cz7ooXX+4zjsl+PzWX9f
k1CUNVW9WKrY2HTvOxQBkGzCCay6J2KxDHG8Xee7OzMuHE+OT5u1DyMVGB8MV5tclvc23Kt0ghQ7
gpSCdrw+R/fQ8el/UWKpSLy0G4GCH5Mlkr5TDy4FU4SanGPHo7urs3kcLM51V5IT9Bwt+Z+nRm0x
sMWS+r+tb4OUbXgew/E1nsyVel1k01VFs3oagVAB2aGNEG0j2bxx1kUxOANp/LPcek5g+9RC9ra8
Z0sDdypvpkKu4PRJqRW1kdW29OYZlYSOz5Tb7VxxBWCz2Bw2WjPG7y/KOPnVBjOIJQKKoFzkRGs/
jaw8ufFjNP5fxE2fmiK/e7tivTzabzK/6aLNaycbkZ5a1HSIWNe0OuXmp/cZo/wi3aZMAdF/sApC
uRD5Bq02hc/E+wyMbBlnJy5WCqTj5xIiuOLLf84AXG8SV3iX4IZ+KyTHzT2kuj2ZxGOreZ7IeQAC
6e0LU5O0kJ/wiBhgWiEkuHceV0K9T/N2k1Lz6NhpJmuGOYMGg66SSVOXVR0BQW3Ppn6jFNFQQimN
GL6WOG5ioHpyrtWt4EXxqz4sh7CxOCjwudqUG0atWEZncKp+uaWTz3R6UTA4PVaqhxvBuoVDMJt3
VM6Ech+MWx+aQZ+8tfcB4QzLfKDDlvXSXAsRRWMa0dQ9WrMRwJrJDMD6jrITxAA0r2mHrrXAnuvV
FcHpDeVxc/5KgwsiKbqwbEsIIFycnKjDaQ2tNxiaUQjt7XWBF+eRkcquIvwhDrv9AcG+vaQlQLoM
TuJCe38EH0VZcVcaMtKb3V7xMga37DvnVhHSo4CfVPka2zCCOUYJGjLyxVPkG/XeoUoFHW5uPtAA
SDfFVrhHKNDbR3p9UauWFRVbF0WGJTGXrijripUS/F7zwiJngw8gAA9AtGGvcWYevpvw7hCsyzoe
uLkDLG4siHyx2QGEqGXq5ziK2w7NVTJmqlqmrlXgc9AoDPJY2x3Hui/mI/tj/Ds88rToVX5AxTrA
8pHV/i5TrO6lFuhxkJOQaqu1dVMHEx1YL6ThzqrLscnn0+jYhOGXXRjXkRB0/VDjEfv4wTnmY7yB
HdNmwmdiE5wvw/+DdxaYUAGX/yiWwrHS/tPuC2QdrGrWnGDR9mKb//Bxa1KaXW3smPTAzvoEd69G
8ia9p9AQSXgYti62PZ8tTUFCpmnLzTdLvdNRKDF0qPvLvMiofgLpkQ3o50E8SXR647lo9RwMDPOL
we2687kNJ9t4sm9UwOkyGFomBSWE95LaSuojhloUZ6z5YQyIiNhTmHECHiXnC4KZXhK7O+tlkVNS
6+7AHj58/kNP3MKadv33ZSKeITqfpn1Lutyu2nT0R28alntTyIIQjgr3Scd+NiG4Kruh1LXkgQq3
E4PZ85tzWQtWS9azJlFwrWDhA4+SFxA7qQ+dWdBKtn47dqWRQ65D1zF+a1Zup1qUPNBdO51M9SY0
ziRvu5DC07i+3b5mke/pzFBjY36c1OmxgAvWIY5VLREnB0c6+c5aMa8eS5S7qX1jWxng+s5aBwH5
UnyintKwm8R+uO6fdglW3fhEeQCvinQB6VsJTYuycqguZ5YW47Bzz1Q9HYR1A2JvB1UF7gXvOcKq
7i5TMaQ9piMpC/5G7LqQ+phk1e4ib7HmnLT79Ae68jm8jZF2g+k4/elAFn3h36A/pNeI5mSF6fD/
b/1RANIL6fLGzWudHC2gj8NSoM5Q+FuUJoorxaLL/KlNCUf63wN9RpVvZqDpVH4e7/2wRWILIvSp
5QE5s9bIsMpxmNns9c+NgpeBgrveAJGBCoHXNc3c16pUGXqt/Pn47e7D6gBJ12eqyha9Xr1kFESS
H6eEL0sLRnXsyadrNpW2KNNe28R3h+SxgLz+9Teaj0yYJyNBh5Ew5In3NTRLkORbDa52L3Y3yiUd
Ox8kBf7uxQFs5T+6Dpv40c/BsWhT2BCc3n1gBm0FbuMxbCNwmuNb7XEkVIrTOn9NKsKpl+4e7uVz
tky1farnlA8wCucFy8uuhL0d+SLkv5YFtnqh9lQcwuTee3ewXdKL5hxGXHowjOgXF4i7e3xe4Wmk
A3yJqiBwyufrZGRQxWAYV43tHIWIFO/uc/rtk8EocdOBGmH0Rf2m77OirxWPzdpuoT8buiyD+wly
SU3kSTXXtOl9nTCNfzgCQkk05017ReT16xx66v60d+9enJg8+7Vi928H89cmg6HQ3wPJFeb/Oqwd
mHRAvv4d8X+aaSz22VqWoE4ObIoXNoleYG8DOEvB0zqohNfbCAWU3Ax39QWhaaLctXh/+B4lvHom
3Izf34cNnkqhQ9E5T3L2Aek1zf4TJrbKGm2PfPrImKByGPxxS3B9bbasxm65IUYA1Po6BUikwrSQ
EoGnYVwz79zMuXBL8IyNg4meosgKSI7hfzlDfaElDU51q9GuYPvIq4/VpiMcpl85BqKBjCiQaHu0
pDcrrHSwAqSzzCSzu0ei51duiZ4nLqIuXgb6NZ+Kw2TINbnkYId02Kd66hNo4zgIDbI3bP4wsc8P
+nigzcSpBLN0aHPSVE/IEb3zoKrepqzAAJ3LEMtwkegKJQjdtCBbhCjszBkme0/EQF4spRbRqXMv
cM8t0x+V+zNuO9/zU+rzMWosbw3UjjluxBj1Qh7RHL9iRqiFeJzFYBXCsmcDCXZCPDfAeHJMqQKF
BBbVQ0BZs7bQ9oZrMOguV9rxU9M1LsNHR8MUyRp0ljmU5Yr4KUrzYpKp/2JVfRw8q6xC13eAohyq
KCdf6+5W
`pragma protect end_protected
