`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2023.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nNXXNukKkBkDVj5EIW2wHPvDM0ZakVbrwLp/zyeg51YxGXiODB5osUXSJG2k4zvQkdQPPCzT56jF
nn+v3VSs8GH4ZlxpwIP3k67ONdfU8Snh20rPZX4Kp8cgra8NqRKMzNXnX8EpXuoiHBkZPTzQKYV1
lTFTWKS6ZraHkxmmDXC/GlX4EBG/+OKjqNyiOvm8qnNAV4V7pBZVoq8apyUtZ/5elWMbslniB+vx
YMBlczQvWqCODl+g46imVjPcCO/5TW1MABrDkaf9PVTdaP/CV4aO/ZOgrVSjF9DkVxJeNFTtI5c8
MnFvORRP5beZWwZQiuXq5m3s6B6acCyRP0oB5g==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
h/HjF2s34dL8D/8sfsxhecpUICVGV3tg+E4O/GsjZl3YEED1CHbzD6mu3E38Grkrq4TxQwxSto35
EitZPcM2yWZgFJMgK+52+HJhL6J9smdK2RZMYusp6+ooXNbkbYdj5iaFFQaxp1q6O5DRFFUc68rY
x/Wmx5lEU/CyVrcJJrk8Mw1G6P2ZLXY5YRJ+3z1ni9Nf7MkGqHyNYy7YDRu20P7IDdeASGl4kLip
KYmbemHfSQPKotEm6tIsO2ekPB6OukKMrpVoiJGXOSqYrXzeVxMHLo/97j2Blx/JaN+3ik60sI3z
buBSYmIZAJ00ZA8PNfZQSCdDFAWkIC/AuKYAV793uN4Z1ysyrEsU2m5iYfr381ZxRuxntVKUeu/7
zLsT1hD38L7eDRNC41fAcl6Wtjvvvtysspb9ts6R+LFl4XCh9E9sVIx4VwPzQCfvArjpWQbk0lCy
ADrQJkI0TVfrfmFLcYunqi+EJMJmv3YB20ZRZzDNErr28+dWAXZfzs7PC5m7MnrjW6VOyQFvX6BV
J2DOMpIPsug1aA7layJEOB04B3ud9qD+/5v25n2R9uYFpVPOvlMdHmVWsS0jgciY0/nI13VWaPS8
se+WOdUkTGwQOA3u+/AF/Fg1/IBf7F0MeItatS6u+jm5s/kyjhGt8B+/hoXWx88vpN5BYKuts73c
YfCMJ97A8XjryNE3fgTwKOjAcbB2+W0HYSqMFRoM70Z1Pk9XANWKbiPejGtoP+z/XIPwAaVpgIua
OgcjhHWvjDEUShFcJAv9lj03vqVJl88XCHv7lSctzeplCbxGc2tfBEjodjZ0g3GgmJyk8cdE5YuA
eXNW1ybuOcVHiL4mnU7IxVVifuORjm8RwgwR+Wc7B+aA2c4YPkksTnVXu2BRPmp+vkhT0TIyfaWb
aOfLliZda9Av5wKpa9prgJgl+O07aQ3ajgyTHSCKKPZ4+XZuhIyCF2dcEt+YweFhjtROw8UqVA2R
oSI14uU2vtaX5E9SMPVsh4rytsHvowKz2uZqmhR1J2k7RyDCusaCbriIjU+myCZo9MGTegbmFiOl
Ii0GOrafTim3JdvkiFMkU0uG8vT8js6OSbPvB8WBDH8vttSAenBTPSu5786hsUSjxvhaoSzZ4h1e
8vkzsBLxMD/w84fG0uSSA3mp/Khel8QKyjehUeJQXc/gC+MKTEQkNY0DubIcZjJQWSDtnAe+Kc/T
yfp3sCYykSlcoFEzwJFIYU/ExRtPc53RTBrRaGuVwcerIt7WR4wfc7CaPV0S7q5oAiIvnrfJUwy+
zECVa9NuVBFvFQq2KpI7C5h2xezQLiwKDzhsYZuikxJIHE2GHH6Ewk3rT+CnykZn7zAOlaOYeXIo
kFVoRPYKSDUIKYqIxPUURBPuqw8d0HjaU/XWbQt5TjQgqq+EeOLwB6bLPNniEWGStiqflKsGY+G4
YpQ5SVGRxqhld2pVfQ//rowpbmoogD8WDyNVgZCm1C69WQtlmVkADbMH5xIqWKt7oa+PfNjoNE3L
yPu4c+sfstLDwWj3CyvywQbJAKc3GhrD6jvCCeVlcPBdmDI8H8btvV6FOUW9atIXJNvmhcxqIsXb
RP6J/vcylaHzrRQ1CQNghgv5zVbbR3GtMezKjiWOYmiX8PQZp0LVGArXz5ECgR1a/Xyq+anpQqG/
sdPs7jlubThoCPg8mccxlB10GnPvI3EBdI8lMSvTtnJMgN7Hf/pHA5mrBE99EtbZsmzdRzt6hGjl
B0F+MvjNpgDIKqRV3VaPS42ChFSMvEOZGYGS+SAIvnADOtSYEdZ82O21/NUgOTEDA2JfdCSBgVmF
1tw8tJpWgM3OEJZN17328nBdC8y3DJSxvG7kNh8fqVDARMPh5Kx/RyVDqit4JXFSZ9gCWgmvVALf
C8dJ9DU0+8tIQYQynkOJW/tduwdCZlIJECSsQTnKj/FlZOyMyXPwSfHH/5HqQpPCtS1osAM+qI+J
0SVkdQieIlHlziNZR9JzJpyTg1DoSwtxd4u11B0mpOn14vj0OX5sWZ7lNDUk95ACvIedlTcAUd33
KO6tGbI+vUjiG0CzizjJSjhb4Kuqmo00bb0lnOrvV9THy0gvBGdtqo9wMk06S6Quyi6CjE/GyEVG
GYs21R3D9lgNBQ2Z3L/eSCjUjNGNWZf1jqf+aZy6k06BM/LVL79hsVwKwepTuozJ+r3Ubye6sRBS
EAFXVAnop5rSTVEIxxEayFS2ldr2Cjo+aUXxZLyQl5JHqLiFqA4CID4ngn20+nIbh/WeS94rYPps
4ZiymXZwjQ4PWIlCmEqnjQorajYXjukqGKDwGJIAwKnkaH1O747YJ8bOqZFFVGBYCbqwFhgeJeVX
XviMuP6E/2KRcAHmm0bS1UEZqgsuYAlsMD2QVoQVg30uK/uOkb0xCR8OPhNoSdEkakomoexNlefE
IQ7DLduXUywRp/Dbjv4Xp6Klys0j5vP+oIo4kAd83KimPOCv8+WahqB+RQ9AY7HBm2cRP/gdiKot
gTYcEYln62xHhvdqtkXsyduLrRFblbKjYxjMyj5roMWrOSawhQVgpUJcry/7BxVphzvyyZzkLLRH
2fNi2IzK9AArCgCKl9dmFzDUJpJtPp2vDykpEN/Sdu6F9TYtzO1sgD6WxTa1GxP0wQs2Oxxro2ar
O8RB5TfoUrJlREveK3d3nEo9BX9nIBEfjQeJ03l9BqIviUtqDzdmapFAOx/G4xbiNFnac1vEZZTx
DoSzg2E0tkuBw4ZFv4YIEetKY0Wte6ZsnK0CxQAHvgqGzpvOX3PGcVFKMHctbpgkzjmDf9SC2r6w
URmxyOKb3nmrJZA3Hp4kAc2kLr9mjxBoqvAt+s9ZftFQeM6yEh665DQ8tRbuGVRzeuIZEZTg2nlt
OWqRoU6MDg6wQsFzl/8v6tE5ZbERAV7ccWOyCEaklVv9NNWdod/c11ilSQa2hAEHw6dNdbzMlGvZ
fflnlJ2hzZHhxHgrfNA2Ldwzed0tEPlUTHHYCu6pHeJVPFClr0kLjxDahM59ZDWeBardoAgGR+xn
zj2PRByA3qpg/QMhk5B1m1LKp/9J7qcyv7dTg3uiPNJHdRkkjqBQZsrq3pYElyPSmSx7HH74L0LG
27mGl/+WgJOd5T2tPHJ/rNKMSgv2nnfF+m7GeMmr34Se7gyr+JKkOZwsoLXlA4E2jTY1O9GQJTCP
ZlzVCiq2UbVbNHsJpXl0VCVi9Snusq+ZpuxMGr4BBdjvnzqBihAu22SdcxxIx2MXXkhR8plVJgIV
DC9GacKIEeZoq7v9xj6Or24FKd7206IoqfusT2j57KSKHsER9MZzpGuWytf0iP+iUGUXFdLZiksc
kW2Ld8LER78l5LRqIhoc/Ij2XKHW7/lYmca4ZAhlQyNekrR60VBShytU7b6f7DA1OUISmTixuOce
8+5mBBPNIxmemPoMoP3xEzrbd6sYr/PSytH0h72sEUt5nqqVWYBYJWkeOoOhSii+PaccTUoN7tTd
PtZoT9tNGAXH8DCShoLFWVSlRXBL92hViFxYmgpRodmOg9oVkv7+PZix+raQi8UCdxZM/1qZ8Ae+
qf/1teCJNCTFyF5z1z9aYWpT6W3uXKJPQpRNlFa6sMhbo+Qv/oYBV+7ivdi1unnFKPxQtvPDcqJg
NbpNbKH7P8CUJZQa1zj/WIH8oU9Gt2ImouyxA1iQSszsu3nsebPxuMWOdk5XNSZoTAkaLrBhKHoq
y5Rb+ELOVcBhheLx3AohVnApbTGXYkhf9ELBiSTpfJtQ5bU6Wiy+opmHRc+1oGSLxJZsmJ3pvXP4
ys4rB0DXnsRWuWMcqM9olpvUKUWsvwJzLMV4B51xkIePuaBXA+pi1X6n2EUwtm0CRInKCYnSoywp
UII7+gkM6uvEnNfIbNd0iaFsmETCHb3JuBP+KB0BYiOX2MdcpjRs7CJrLVAkqJYtOmc4khQJiHja
nRSOmj+b1oCPNb3FHUUjxdi/xywJ7yGles1nobNJI1Y1kZ5AenZaQn4H8GEYzP8pkpUFf64fyL52
Qt3Xnz4U/8kTHpxZFBpRn6Kt8euAtM1mcRDg77v9Iqt36yaYyNmPazHGWGeNbEOe8t5cWfTGemaN
1iFjM0TeWYC+ndPcyLKYqcNo7OvTFZ8SjfeaRsNo+Zk+c0Wm945rg3dOcoOMBXBpp7mtKXV/Ajh5
fmeAcfjWUysG1DhoSOxEHy/sNdmFYsufl6ywr+CVHYfYtW07XtwbQ83aSWP++h6opn7qGUjqSB/U
pY8dlFe1ucL+6GXXVwhIRNx/y55MjQ28AopZelG4ozetzHVhZ4FzZwwQXQEDeB7UwMbGlHUxO/H4
gAxaoSLv95kjIk46hbvMD+w/5+sCLtGTImaUcjZZWrF7QvfRhphl1jpwNrpzwGO6bM1i/XoFFcqQ
bSCuN4GCvr2jMoDQ5w+SwqhMczDr7uWwWjCEr0FVbxK4HzpCNTML/vjiqQoztu7nFGf1c5CMJ/+9
UOlCQUwD2YP+RvsJmesuvv7kpmqeVZxgnok3CdHlDPE8t3eIMKjOkQ6y8dVKA8pXLljbFPB98/mg
hnS2kZUky1jGJwY811gNVO1cz8pgWoyuPgtmK8bWgD0szAs/A+MT4BzwG8QLmLQosL2PTuaF9mNU
MTDrrY4fghfrXb/XzY/5fswOH7ne9aHUWQdiq5chh5aTz92Eanv2CEMjn0Sn6XAXtUzNNwlklQ5+
xiHxtnbc/j67KhAL0eIsCAEPWFE2sHl6Q0849To7YnbRoM/1dRYpCnRAfhEb40rOAzfTOMF7HuST
NpiQ0VdnMYJ6mgrxqTUKjXHrXorhvbsTvb/KsVPxsgJKrVYj7jTf5usCjgMDtT0BNk+8sUk2w0AF
qKXs/+Sjd1pucHXpJLhllCQLUnN6NGjmeUNeHRPynYO4GcU993TR2z0HLGdPL6FWf0uOCO+AXsYc
yDkH+XdpZjI59HeT8bqvcDSaKIY73D4PLIE6XwZMbmlHkYZ5OOug62LKAXixt/zdvQzugOntXvhk
khd19jBZZnS4wFMb4imNxkSWjFl4yI9rK81w6f7ufIhbDA3dZVawwNDW30nrku/XOvY359OPgyO3
pumKCyIyVvzC648GfuU3RhjqgM65LwJBDH6GLaySHLDwCb+qe9bcSagTvfBc3jnveZyKccXkh4pd
rSg0R/dBvnwdBGRT3NYtycg8Q75lJytzgDZoudR/LMmQPFrXWKOl7czHab3FrVVGM4m5p7BH0LCg
Q24kpwDS1NRRdHVf3zpidFxjEFOz71sHuv1FWikfB42NfeLjNUcKcLNbXGfPaf/tcrTOR6kafA14
o2H+YsKmWO+CK2vc4dfhpdkAZxY0/HYIOC8mayiVPjt7RWy+ud8gtsmThViECn17s2BozWfMwTiu
JlAPRYjQiUvt/ck+Qxlb3BAEv+p954UJHeS6V5BPzBTHterI1YrQYg8LSTJ7JchaxKv8imTbywfD
CieQL6+cjVQd6bGQLSZyQ09sE0jkBIfp0TK01yPyzyjep214FLaMbhE7NBZjUcCyperuHFfco2zz
cwfJ8phloDr+5LSdnKAV8SIMTLJM5haclTekItRpYmQkYUDkgG/yvnj188K9kHMvdAkQK+YsDBg9
0eURyQQWzOJhl9wqe/F3hhNUizTzqd8RJ9zafEW25/u28rhcXWlWIGQdVcb7wVzO/LHi54JbNObE
R+POroKSSQ8gnlA0nyuxKmQ9RU9MH3kwP15G/J7poQH9rEYknVRjchaIK9UCF4kGIHeZWQVpojv7
1Xk8zAmq17AIyNYxPSaQQzgkfbQ9BVKZ9phVfmoah/Aw8fjCDGwkgZ1Ck2buAbI/gkF2mgOCcq+z
wEArqLmLdyGcjmTn6edpDebIPgwq0oGL6KXP6vQ43dEA1ry1nlUFOdLHAXxwlzQy+TnQtB8FxsL1
NcFrznFLNjye+LZiOVJsYWNA+x1c/auvRiaGEr0xW/nXfa+1E9GEr4KrmyhLaWdQwHLfXQf7HdHo
sMr0/vARcVS/+UR076NiKbV/V80g1mwkCypwoQT8Joa7wMDTgcrM1RwBkptbTwfXd3Z4NS537OAx
y0PmXl5x3tpOFugbU+UyPyT3PzxbFuDZQNndHSSxySEoRUbPHUi4XI/C6q4akcp3JxazlqXDv30s
6Fb5XrXf2JWxuIlNQWRUF9LjQHogelnK8oej0/3/RyJKMFQrala1vaZpVtH3r/RuRXLJmt3LyyOW
XYxVeNVqi0orxcNPioJonDbDYIGB/5aWwTzJt2Yh4e+6Xqr1z5tQltCRjkMCkf6hRAQwCOgxC4Xk
IfUGESN0rkc+qOVT5m2lBH2oopHc49C5e5smQSeHL9QkfdqMvW2B1UCyzoHCEdQRTEI4i9V1vnlf
VRFiy6ZsyVqhOVRt4AqXHn5n6yTNu+O2sCIpO8S7aVYvNXykofeVldY2UYRJGvgQK5LoSpdVxPIb
F/DIIypw3tCGhamyQf6HjIXAAunVx2cEkJ2ULfP9ixff/xzLRBF70OmKFxJWMa4IwBktU38RG9ec
CkSC1Q/18QTJ23KOFAsVJJ/98FWpjoqcrLuefESUpT7ZiHss9NsT7QN+K7MQx72z+JVq6dWTUe50
RXMP/itzYH3oZ40FicjOdOn0gPi8/67MqLxT8vWaUkcYoAGUVS7+ClIKc8Jh8jrrKIxIxDPe9j45
ZFZnfObwvy6QmdcY9kpLPNNfJU3dI79gTaOduz95mx1xndx/Xtck7CoHHiw0yP7JzhIa32qFl5gM
n7Z+mIfR+xjnzUcYaxo47bBVcq1ixc07pWZdHuH+8jNLElWxRyCBm5BNOi5ybA2pdRMEqR/tksmG
YsvKtuFeF+mG0ZJFF3CurffEMrKj3pIW9v1vjJjpZ0lBSlBPIyeu5ralmOj82LDGRJWslFm8TFOq
HhyX9CognJdFz0NF0Z+TouezVXKDutsZqgRbiHxPL3wy3nbWHJNM8UeeD9KN7ILrpzeyl9L6DUUC
PSVF1Iwka7wxGYA4XiA8ipmzpSC5uyP3z+F5KYtZM1xgPJhZlzilj9Kx1/GSmixfckNZSPTfLs7/
+mhUfbZQmDbybvBZu1q+dzit8Pi2ySb9vEsN8WFt4MbOUiJihEr4kMk9KW1RaPkNNrsSkggIKM72
ljqS1gjmqUgrOiH8xMlQmA0oxs01p3HqDwewUiYrRA4Ge4qpk7huw81N7J0shq4qzdoNmqXqkplE
L48xQd2aVlaFLVldbeh/lkVjsKEw/NiCtDdUHZZJjNSLFRROHTyYDnR3ePjl4RI34DEVJfzIY/Ze
TkhaUO/gOWS4YB7tqYr4gOQFaOUUVYS2ZRUQ3NXLBfPpmzK9xzDxl2T9UtvBxQyn+SJivQfMyfah
jF5Y0DkNfPZYDv11TFEOZoeN6WfuTU6/pmvpCeo2QtrKWMky5qbtiuwA1RgcR9HP4/NUGAQdlVpp
nTehJ43xoanJyvHwud7MzkUH+r872izylgE5rb5k69LQ9kthTBGvPRXyPMKbrSJvUpQ6gks3Q92s
BAYy6ma5Velo4CDZNnRHcL6bZwyCuh4oUvKl/Rid18PAFpesTUnS47WnYLoYbgvjZb1l58QFF0E2
vmHsoBOj61Icj8wOO61M5yML+PoDMDooEyLxDNHU3ARl2qVctpRTv5BhWyspq3sAnWGb+CQqmJer
FbZc0gbN7xZRqxU0ef+Nvl4xVKg4PPCUfb1rlnbMvGucGFZfySqXIw9j8AWWcr8IcqGseduz6pSs
FgLJLV7ry0zWSA3m16rXZxNHtfiikmkMhiHLZxRgcqaS0dapza+5gklur/XkR42QCNZElxLp92tM
YVRA7ghvcnLyXLrZ/p9ixboeBmbEg6ncQhHcFmmMEyRGhcfxrDcimvLsw1LItoDqxAKiV+mk+NV8
YVONnSR8o7dHUMeaaa60Ji5b2WKenClSW5o+nwtLK96+pWhZExJRxooa79hGqKPNUG5OYVOLmwPd
LOP58W8VQTOQ2yud0xd2zDhKbNIX3vNRq77Feh6eEoKigZb71IHLvvHjvggwfVtj529IHyhYN0by
LjqWi/tzqC31WJ1l2me+2JS5IP6/tFUymYBfMSDDqhuRA6pJpY22oV/Elyjj4dUxQNvufcQWk0Yv
X/Dj0NfzJAaanM85dNVp03xsiYsqq3pmBPXysuGKTqU5RSQZx0PdiyVHlN0hd1zKAJ1ioNoQRElj
JeaGq8DyWTqB+LBXuDyzAHRQ28NFErKd83FrK8QLZhv4i/WwoFuddwmMhCp0FPtU42JIwrJCYf+V
z7i2G4/c5mifonS6LBAGcrUCdhGZnNp4NJeFsHgX+en0CL4jeuHyiAMsDtjhLQLzb3QwMVW/yfyC
NTzoY2JJ9mbpmnxG+5u2Od0Qx1Ae5lXHVMktq0t/iU9T2anM5fjwN1UFLf8oboycPyLgHEwo4vbI
dsjUFVF2dOH0GmMOcfJSS+Bufj4jDFu5207fw+4VK3kIZ41PFPZjgTvCTiRAPaHQvTDiBfO9WW6A
wARpVqo72cElmpogMx2X4NQzwdGOs7bZgzWVga9fjzzTGqr5ZXD67Be+fH1Y32l083bCgGbjYHTD
QXo5jJ+1nopVkkFA/h3FJ1fltQJyJW+SXhZmxM4CWP9szcBO6D3VfC9G2uKsP1M9dJ6WjLJxBCh5
A9r0Z6uxVKSYZvEHjfkR2eekyUqhRczWsjNeI1SKINavT1/l1Hy9FStHN9SYpSMX8BCbULEkgTln
EAr96P0Gnzea0E6CWd++m3hY573ivm/hJRdDyJdzMicZV+rRKoOe/ZT6GU81kLp44k5ENkXws66M
6VT0UcbllNq0KEGoNKqclQg+cERu+n/Or0XEsM9wo8r5eMkHkDVGK1FBbitQhqT8Bv96+rpLEjiN
5FLKNA5g6+yBFQDgX6DKZg/yab0aWyC+89j/Br8NAeNe74qdOdkGlx9M64VeWN/Fl10Vhbv4FSp9
Kvb4rs83O4xXt5rNNWOu0/I+bzBiEjw0ysZ7awZ+v3T4ZfQENIQRSY2lMbgbvvUgKJ/TkfWRpYZw
2ScolMJYr2jTgK1gjnsR5IKWRdOyOSyxs94VebChDVwJxz75lruBtHH1VpGKPc1u7K9WuKTDHbUX
EDH1vTZnGNejTV96zWad/jRQkwe+8qWkiAgEfNPCWEy5gtK9FSCYCdbIRTLC5C7nFrWsnqIO6IU+
2zEqYAwMeI3/wpGR0gUW2oyvSRCudn3UpqbS0/8tDm1NVcSp1nfZiGHItXyXKFHY4szZC9N3HXTx
e3Q3buHTzEpO1GM66N1/TRSWWDrVO+Du0zbB3uoxL4/ySuEhxu2b0yYCXgiwxe5acfwLge12xszQ
wQ686XjfJ2G1T99lChnOFuMwZaWch0xCy9uhQh0d+KnrWlsEKg4YagIicLOJJLKvjzLSNb2sbTVk
7zr10Rxt7mc2nqVY81qn/JAKeMV0LtMrPID5xrBWo7MsBF9zmxKDH3gdx5OH3DUjvZKIPL8Q1cTV
8fZ0amLhCjSFQqwkVoaRM4wPkXhFKyT1+Dd6quFq1+QzWRvpuWEr/d19P9tsdZji5XX1flHu04bG
ZSXSkXt6jnyBQIQwTdpV65EfNyqwgdUXkyoDzuIhvKAabxBE3az4XLJPCR9O5MxZplhp+0zZ02C6
BA5mmEYsxxlvZMnEzxlq09el9WtCMb2+0C5MvmecKUgU3Ne0nV7BCATmn5eduN4GNFN2Z0QD7Skj
EGp5PvL3R4QB85KghgC+MkafOC3BsRpwxuAAB9LoSh/IfjwBs5LM1vTQsz5FrGObxuIZmnSIGmZV
34hvpCoSMGePHgK5SEpKFL3Bt2YazuOp0msXCD8xuue1Z+dNIU6/2RNbOF2Oc73zM1XXjByXUSNY
M76r4pW2f5UKpk/i8/oiiUXD2QCiNofdFnyHb0XAG2hUYPaMFWwHRkeyn9q/6plvgJTA5E3hBH0K
0qOzLCB5Wk2jS29r6i8zdO9466PBPmiV/xMwZD2Bf8icAyg+rbyPUD38QDbNMhVJQts+Sm6nKHGJ
jy88e6JI1qTyLtTVse6UPzB3TVqXKbEF+Wf4alIHm4OPk5hmjiIsYqm4asEj20gPrKLPdcvvWPJY
srykNh1hmYyNZP1PaMDVrzZdzo1D69j4ONhM1CBnVLzSdY+7ZA8y+FEFRXoXhtz5H0Ne8LfxUso6
GD1usri4Ag0LBaiuMXs+c2juUf/Jm1g8ob1ZgYiaW0kkORfD2cuhw+JWzQDZ/CGh/I8qQvFkkaW2
Z6MGa5+Av7Hc7XwHyo1UrJa868tLojnoXnTqfMcrA7HlFugRVVoVL2A0C04BcM56WuOD96L3hYMF
FrVt3X9xm8rPkOC/8672Km0rM6p98e6LtRxNl5lCRD0yTW1eqw1JIMeg3X4mOyyg7kAnUXM2MbM9
u9uqrtOPP+WjfLnVpKmqHkR1KVvnlZ7Silr9B0zFDSiiP9NI2J59idNF70Sn2wQzykVpDPpvmq5O
VdBDJZ7UWgI1fdVpMhiyo/OscIYyh4IuMYS78DoTIpG3C7hn+1unBm0rNKr6BqNVC72qt241QHzl
zujw5Uac9uKI5jkzRTvu9huH20bGf0R1V01zQ40vORrCvUnn6KOvb3zl9EGsHhLFUPbAVuc3GgaX
AlPcFozWOIYau2egK5EvvsJlygzq/20Ey5IgHNIi7BcrwFK18Rdtd5YgZHZjvSTL0mEsPUbHM9Mw
wJBlgq3Jg18oyAgGs14Qkyj6jDtPDYjvstoPgPRQCotA+mcV/KfjNvc0av4MLmYXhgTQbW+hMkBS
vlTuMwLOvmGLJ300kZk1cqGJ+m3/NscBpn6d0uJ5DPKb0reTy30dYMrvzsm0pw0t8kpP2RTFGhQq
J+23qmN7UwxkhICvp5XEgFJs4stllzRS+hrzGWgCZ5nVMnqBDmqBuYmvzBuqyIW7y2EBYhD4XbpD
L3KKCdHF4snG3n6jkZ1hLn/ktO7Fik4MxO0Np3Xb0yI2RAHAvno6EgcBlf1eeQxyN8fmtlYrrl4C
sFSVo6GIXn6bgADt0RjPoLW9WxvjDr1zUO9lBpbRBVqNLm4cWbitJQ2DQc/CYHDTzb3hZyrDES5/
UDb+ekRd6Z86/H7HAkJ7l1hyAB3ghACoEQVCPyONvsHUbbAWAuIVbJ70jEYqkvr4RcqhCg51/FRL
Hnmvx90y9G11AcDXMA4vk6jN7CprWK1Z19npjHa2O1ZnJl2ih/pcQxWoBkI7YAeY4t2GMOPx3xUf
No9ZxtrNqRxdoHJTH09DeJr50RYYdnJGwPcpoymmWcOrGhQwPPTH7v+0FijJH2GVfs7O+OgidkI4
NXM4DYm+EjB56iQj9wuvrzR9aHguk1MT5HnwDKJLDb9gbqfjFPeY94pP5JkRcGKy+UzNYClcDpzJ
OM+DT83KUbI/AsTVdcVQDZ3mfgMcoi+BQEFMJ3beE9wddq1ar/phFwT3ZYTBLyj/oWKOpoWS2Iap
PieC/RkYL+LL4upshUzNmlHQwAethTxtXCWKhOX7RpENt6knJWeGYeniSfthDSh9kKcmmbHuZJNm
Ea3kW34srnDUp45mK3f8+3pBDCjFHaw8slZhMZOTqOBmSaDLMhkksl+heZKC6HRe7HrFVuzDzNOu
X/nUgB35nhUGtexgGgdUtfI7FAfBNJTsSzibY5G4dAJzXeWDIS8UPjy0y6z6NqbECAsxcGg6J84p
WHmR+l5r2GPNU8jcIzAF85KnwKP6pV0e5aeW40su2QkYkLjjxPD2hO8Jln7idyYcIfW6WCzcGQ3J
N9LPzGIU1+QsyVhkaXgqY5w4WkeLw1HzMHcKfrrqcHyR9Um8D9M74DG2jNJVh0JDlDIbyyZYjQsV
3T++zidmJ4uIZDFlvsie+AE6QKNy62bM/bD3r+jd3WYNAYUhFp0ZCnomGHtWQTuqFd4ppAyg+UzR
cmNNwtrt/gyvva4obYjiX2d71nVE7U78CGzLkwM8YI9WJqphk1FHbBsPJXcKp2pN+hDEpxl51l5/
SCb9rMZTIuvjnCjMYdi1m5UN+GEeA0R2Wx1VzhYAclJxXI1armXnzmgWG3Waucuaa4AYQsd60jDM
TBvmQYBQxhyJdcunjOm6lsTlwDJaVwI0ucshiv6lu1MWoPgt+p4WFEdqGz3UXjhLtcUVptMkWAxK
lAW8jNBt6Ro/dCwoAI/7dWykQ4zLDUFM9bSJugfgDHgmRPmhXnu2gj5/zFdUev3s/1TtyeO9Bdto
b1JRrdg4zjCJF1T+r3omSQDZhpmlIqGUZ3p8v64KYN8aSocUNPhkFb46jEahobtw0OeWwvFmhQo8
tr5qX81uN9BuDVh09rn7DED2rmhGO2hGCyh9uivMAND/r4vJygiRcD5ym49Tas4iocYTrMZOXNoP
hWLWy4HVUKSTi5c/GfVtW3GIP5Z5o2NV9ROwNB3Iejqq5jmwgRjVN6KuKKjlgsMXvJMKhRYzSwob
GDfnLhbHUKcZgYzmAD0MWOqoYfYL7CoBuWLmJOQ774mJh4QP4wkiFnesnn7ZHrKIWXWhB0Zkb/gk
nI35VvKR7XjthHWoQ2nt714sAiI+LlzXy1EKYQEbCstXNJHrLDsGkQqPnbm7vvs0c7Sg14Sl9g09
F/ny/R9HwQaUCcs5Z9GPO1LmbciDKLwLe0qxCTYdNnX5czpG+zFM5IM5yXOWacfTW92Jqw01BedT
OqTNpQHO3iDXoJaa58Df8Uv0O3B26U+I5tc7M73uwOXR+yNnQYIhSZY30VtmpGFVV3dGf7XFAFxw
IvycA606wiE1h0mjCYpDWVa4KtfVtZB4M6Ulrbdgu/dmn8CD5D8MDmVGqeMGBJ3czYi+O9Whs3+v
Uz0BIjGAu/8wk8PTsK1zdYgU7d4qpke0GxWejYEasUluL5THI3FDoRFb00gV6LIEmCgsG8UI3LzU
jSECT5jXz/syKLxonC28L+1e8XcWthTtrURxHHa4IO+o/n+MzFU/8ee3Homv94IgpFt9Ce1n0XxC
D/oer8D5OB9xy/CVE+C8F4lIc3hsWtVvG4kDHzuQFqItGCg+5sxpZ2S3oAHrVQnwCCvRQul2/3nT
tw8xO+pcKU93poTrzgO3FIgV8Xv7RHUNPPOaB37JhNBoWegPNbbLaIjsXTFe9fo3cYvBCiH/YJK7
smdycFePGwoNB05aNrpnYRcyID6+xkVlQjmmZjqb8NNxyFNOaSSWwm5fN033D5ZZr+VNZmR/s8c3
xhP5VZC3u4AFhu3WSR5g+yvkyrWZ9VrNJd4KfNQ56zby/wJ9avlqq8dtjZXWdghxXA5sGYk6H7h2
0Z0eWa93ET3WreJlchBvK90KCG3jSl5WJevzppzEJubaWP2NKjZ5gRLhsVVyIF/lPHqUbBt9X7uQ
rEUIIiRy66qYmlcqBlIOy2Y0gG3PPtcIt8iuHjjd/O79i8Pufg8gCkzRCz0Vy/g04FfsmdsRAON6
f4Sbcg+k1/lPnV1AwGymHfBrNUzNSPlHIfBKcvVZQaDRSh2S9XLYOYHMdBJtEdTEnGKXROnF0R0X
6hGVbPUAH34uk0m/0TmPwr0FmSJfAPyavAu3TuM3Dd2/xu5rgi6gWi/esgqsRF+4PdPBE+TsUshU
b9NPUO45UPjtYgr7X399aKLqVzhHhdjvEKhCRBIYoJZHZAFwb3VQB3/byNGwGUrnf1MjBivlIgJa
cOWzlyWiW+Isz7UgqBdLg2b5t1kHAA0QHUHduyE4X2T2rPiYba4cnX4NT50NyfciLsmzY+/FSXim
DdpRUkNgBtbPw3Hb+OGi6Do3RF2VWWLfEq2yME5hCv/9gOz3tkPqPAONJ/00/loIzyKbigp6Z1VX
Pib0t7AFMzdk58mWnAGixB0pataaT3HV3icZ/SwEizaJ6tJSqmfa8TSN9AKdqehQEVG+OGGNQpVZ
uM5aSCigL5BbiCmLZPE3+ujHQRv++KnJdacHsRbA33LZxn4E7Limdogn1K46C8KceEn5dIEpR+8/
UIbm/InsplNMFhV3g5Rd3B3RMHfYJWgKwpY+4l4Uogs5UnHpaRWh9+ido5EOP8XkyhhuvONAe5UW
0ddxF3/F5TW7yamBJTsJUoNgc6MMIaWVke7hiNWMKPimUIBB6KeFyDXuizzoXk6JVChciGTKKF4o
ZGbpqjkUTZ5IypUtwg4dT7cTozE1yGMaKNHzGV+41Y6bfWDeeDfxFhQFn0o7tZTUKtY8lgAphO1W
p2q1droAKMiEIQx1CU/C6Rr2MbecYAJZHwqXAl+XaKQRsx+OmZ+Dxxbj0M4g2CeQbuYSkC68YsIz
EemXDmVpUnwkdpiGS6AYIqPmBA7BhiBga5JUAGofKPKwHCtVPz4LCX1SnP5AtukGeL0qpW/uMsjH
8HBO0DQblDEj5BZ97azrWD8AAcWopq4QVKuAVrl9S/VwqARrGZKlV0/lNbLGeZXaAB2H3bPVRaeB
AbNWnScvS+Z04zgwPum+HmNxYnButrEBZ9ahzxQOxkYnkT0kk5wH3LHVuEOAc2P+SYmsmgNoycie
1vzLd6UawKlaK55wF0cTgpcKkUaQGk5f8R6wj9lvD0CeSEA/uFABHkTj99NwcTu3BWHsbbANA8rz
kGbkuq5DZhjFkBSfxDR211CbmMDrGsYTJO91x0+OfjGus4KhFSeAfuD6/0JEoatpZhmm+L8BwsEH
J50//La8qQblYVcaO3S/zdx9nsVTLhfWAb6tcCrON8oB4EWPotb7CI1C2zRV9WiftGB4fVPQhbMS
61EM+R4n+RgQUzZ0ZSDVVZDzqw39Ed+Y5u6OfPX6EK2vNlDQZcrENjY6pacAaa0nG4COZiAKidvu
YgRiDg7oZY8D7gHj/VH/HnA3B//nwYwdmDystCz+Y+t7LcGBa36ikbGlhp3IPBrztiNX/Xi/Nvk/
Q3Zm38+LLDn+q5OQpLAFqBx0/qGQoQqjClN0xs8sysQN9SGOECxgxsD2Qg2OJKQyLfhN6Vio6wkg
aEYBOinSfjV09cbRmD/d2sdOJIsNWLQY0P9umZ9IaghXlxHV+THYMC4mP8Pnl/xO1ezB//E8ah5/
Y1jt/hqMdMi6dEljcCdUFWDM5O5+TJZFc28j3C0p05OMX8R6aE4h2aLGeESOqLWx/uYLKM749JdS
KUiOSTyF3tvr9PlE/6Up2IRVohxnPUz7dzv2gyDPQcUqjIx6oit1kYiOhpZ+3AXOxaGZQ+LOWGTW
XH6qiPm4hX7VcBEfb6OwZpSIeQ/SMWLD43RjjMzlR2JDTf1sOrKjoqAX84LU41U1icb5HT7B/7Ta
C29U5tXle+gDEHICehj/WffiWsQvcoTdpMsoqdCGrEkaxWjwg7Wl9GwhKtJY8miIpru6fjk6VYvf
M7jQNM2xsmsch82J0fBtTWywoaND+usjyfLf2Umkj4CFA+Hdf/xzscHsqciTMZeSNIDECIK4x7Gi
Prhvl4L+i9u9hJ/xFO44Xi56LZ3TfXjNQrWrRZAV8YCTel/TZesD8QYELuqW9jVs6fFTamDbAGs9
lJuHBBHQhq/knXImOyIU7LGZpikYjh5n/wPIs23XF/7s5BLXmkwzybSYZ359q4UzwSbReGGiAiFp
jXPoa3cB2lfEmlhOBVGen4S3f0tNb4V9s4NFtje17jIs7xyvbcTqR6NPQfeMy0RXW6cOriQXTACN
FwBWrU5roOGFR+VmkdrIAq+yXPX2/Pbl4T/n2mqxN6WOWIRa2LYDsv1pRCjaGrv2BdOZCnDakRXF
DiDfpcgobftj2t7H211ZWHDArj+fBZ2V8OiP4ILZHqMg9MnhfuI7k9+Fbp3AN9U1uPoZolVeXrXn
M9cqjXdL1Aa3cjkTv5r2ltxCk/nmUx20ZowKhns+t5iSqojl1y5CNQjBu8wvgkCRUWcrcXQPxHZ+
Qbcas9i4csIjE5Ja1mI/xvs1LRSsBMXky789j+AEz76ZlPaJPx2atUsZD8utdACvOEXmHJQJzMzU
4OKSZzlGerjPYjUb5W/eF3Rn+13so1YukchcBf3BWYoIPxp+LkccHW4RoI3lzRwcxhO98MfomIDw
jJhhHmvp8iE1oFR9WklkfCcuhTEEXkC3mWor8PrsnQq5hsCrmP/b3FByB6nWtxor4w1bWcCdYJVV
vNgLwVyA+lkYKRQt7bU8J632AwrEbPJUGvYRCtw7OA1cU+ebbdHTYVEy1pTyg6M0iqYs8QjQT9ZF
6eXNqU8qXJUGiXt8MgRQ/Q6TZwP3eutbXUxT5cBnqRVsheqrP5RnpeO/8c5vC4k/RvG8oXneUeBH
EVjAKOuUFl0UIlq2rbXiXLGy49Xe6O82ibWTbNwveybT5YSe+WQM8VA3N0O5ekozfs7xqh/QwlAL
YTaxv70OMud5o9cU13mQecTMdTNmbqnTmH7xp1AKssncD3QTCFuzLMsocNDz3T22RSowJ1XWogHY
vEsnENrsvrTM+3M6w1/HieUr/culit2DqUb0AA2AN9zQ6xG2wlwkgLDiaJn4wsi40zNKkDSOPgzK
iy41OPoImeN3P8pVvgWPQKZUUTfxypbPew/MF4JlMNtx1Q9UsIyyMroBRhFqDMYclrMmMx9RtsLQ
SzMgA/lNQqAGc9GGFG2wrDrx5LdNkNbEVyjr2nLrNn/khidLtHYDnfbcC/DWZMSbAv7fOJv7YpPE
gz2XiWtn5UeEMIfOpGlGeImmo8gZPan4zLBOdq24i6CejburYd4F3WIpHteIdKRluns9j6gqLJSg
loYnmtJiIb44BdNSaYm049N3pvOKQiQ7FuD4st7m+fqvWGrg6rBUIlJqz96Apo5E7BqWP5bsPaHZ
ybzdxyJGUNVTDmExJqgiTe9HEjvOwFmu51RQIdntesurkPQhXie6qEvhVDRP7bqLdvbDZH/WI7ne
iRam9UvuDfyO+r60pJxyN2pG8VVmpLwONuTShPhfri5SdpfSgwVXlsk0pchez/S3jEuBWonRSUk5
6UY5IKsBYHBoBN13AE47sHDepWDR/JJ8N/I/T5AC49CIZkejXZpndA5BjFsWz0qnoj56HAQGD4Yh
x3D97e9rHcN0aeTzkwJlAA1+Y7SWv6bZbj4vVr7DMIwDqtsxWqUn+JYbnf9ieIX/f8ybAEHnCCI8
YrGKG0WtxZdVBw3esnUo1OV05ekXvHy8dyZviptqbp2x3qJLQEFZW1l9he8mM82ZB8zwbevw3Zup
+TsflU8TmqAtg7a6J2eoZGcH+oKEpwjolYNgE7xpNarhki8/os27LlZNzyBDqoSpzuRhYbuR48i/
/aC16mzJFKhtUEjwUGsajkouNLA2UjQGh+U1WMTIQcUWz31/r0JUcStbxvYdft6CFgHX0j6PAzZL
GfZUWy/or3+QYGrkaS2bkowvBOPvgLLwhAEq73RnVlI1qArUr3YY6LcgCAdcjycmXhyRBRWj8vDp
0DaaNeHOrHG6gRfGNtHV1wUGpJnjeROlP2x8rLh/ObauK5+NdiZmP7MxczRo5//n4E/lACiidvt8
cs5XqmhmIdab2Y6HPzkASHHXNKwen8SendnhD0M0PXd2jmf6MSOyqyGNhBHqWQG5m+OywhWmM5lc
gftB2srTBS/I/MQ/0HQ530hS0MHQA7CvS4XUKVO+KRXUxzf+th4mHILBEb2EyztTq4rx51AZtQeX
vOhdwI0NY3TggNozf2/59VNuA8bgR52W49l53zKNj0HNlmRzaZnPD2yKxCypV+33Nt65d9AfzrFO
1eczqO2k6vfdY5b8i8rKr9xZ5QDLVUG3fHfpCPIDx+uPvPzT+bgCl0OTSYVr9tGyNone1NeN4EPT
AFgAPwnIpiqOQ/HHNE94h7PAEw6MTTQZTNB81BxMVJI8etjrz1hzjvXruzZlyYHmdxfA8EhnAh6p
ATu/VaZxX0wa939pFqBYXQq1Lpk5VEf0zKnWYpmPzM/MmPQRSfd1SrqHojeOoHlErGnN874VLrvk
2cD756IPalV29Mw43inT384I7R5h4T4UAZYlWtdNkzoCo9bTVqYhz/4wHJ6vkKAQjUD0oRXx8d7P
2TIam6Rrc0fAK5LuejWaO6u7/yRmKbgC0YrZWeP3ZbyrD7HqoQV/y5VsB2iV10NKbfBiEwlRpiga
Yg3K7UqhVkxuGwGPUiUItmsn6oFIc/Mtu559qyNOnofSmKwkQHpd6GuYe21WrHVDazkgLC4EJcqK
cu0ipuQmXsmXrwF5zuoTB3aHEiPneMMHwBuLnXfu6ddOuOa66r9GVMFoSq3nUELCuBYZV/9xockr
/KMrh54FFS3/mSq6Kvdf/xij9yAbbWeFHZ8dgHD3dqmWwbzRp0jQkgR5aXIWW6JwkpcoqEGlotDh
Zx/VS6x458ZjImEEaCbMd6otfK+UXdnbstz8QAqpyz8gx75+Ft3LMSx2VpKV1dHbby1DHcczbp0J
cOeKV6IAyNq+rWPQb2oYgmaFPMqUjtGHXuilP0wVHXt76n3g7h8Ggy+foGwmtnKW3ifmFUtwigoD
hJYxteaDJK6itMNWBQA8ydQ/XbrLi+nQWwEEGjF/idxXRusjnhOr98B7q8mySowLcOpEXCJoXWWC
2S26mcJS0kiLizSFT5Oxc/57Mbrc0YCrRfKnlRC5Jz3ij+OhKg83viEl1o3FzYUxDkFz47IdmqO/
+m30N8XZgudrUIz+qkjculi4AtSMSL+jNL8RDQ0R04ezNC9yABBe64982ckuP/1zqeXJ4QK5pB2w
vxT2kwWFl3wobMTY/MouKrxY4L+q65QUcJDzcChHgsIBaGBCjU49FD+V2F1xeZQJHjMvFTc/s9yf
uTcJwZ+QZCpPFkn1AnLVfbDkPrqrQcGhgLBTAmPsQzFz/a1s3ZM1VMxR3SFawADDlpbE/XdM0TnG
TQz+IE9Hc3FdRhd/CTTtuwDwMXkEvplFCXVuDmu5wtU3RatgEuhy+k03YQZbMPHnMQrB1Q7MtuUR
VHVvz2BVm+J2BWoRuOe5zCn96jd7nYqLIdzQQawqdTO7tiF9z+i9NbIujbfhr92c7AwiQ61D9XOF
LJxhWllzaTT2J72wT77Dgnf1fCnSCFLr7uQt9bdx1pS8SMKsP6iifJMN+4o/Iy8LJgV1LOwTJwvO
LbaMihuYMBxwSDfZfOHR4Gdz+Kwa+3ojBPxvjsL/bPlLw2iOwu1UiYNWLkmHPH4p99YJyOX3iqD/
7f+mbVxcYodjmblS+WF/QmAti/SbUcUKXXozTnBadmvz4Loh3ZL7KP7FWG4A9mrYn45KKUb998tV
r3oXyNeD73c9eGfG1xdVVIwHsbVnfmmcAt1lue7+Po8yMXWHa+pBl+r5ZRLKdI09O7weCH9ZAtF3
F1Wapt1d/PU99e3KPbZzMcfc7hOgfJzvQ++YRYQHyqK4UrHcrc+hAahU1Mup/z30++bGUl9w3YDj
MCtaX/s8Y00L0cG5J5HtuvmX83iwcYRdaPgsJA3e5L/rn1H6cjpWkydAa+jIPG8TmMS/Fao29tyi
h/jAMWdVutauYa1+25kqAtFvd0jtNYt5seOlohBZwWwOwpwbM6cAbuXQQZ2EUABtHJMQt9OITExD
x8xnf3fN3qkFiF6eB5uB1/kq0A7K0GKPqwyIgkl6w9YPWKACdJmj48VfuKDqTDx3or2xUDcc+B5e
sNf+5nqSHPfh2mvQM8r9/DLVJIm7owIEFl20bYaNx0P9EKIb/bCfar1j2xoYlXqFKbSXgW0Bzq1j
ARRKkcXkOAK/sqN+/gYrlE27dqAe1U54xmgnLl5lgDswlgf3yM6mAqqQbQ7YgMm8PlciXx7WeT85
h6fHUjysBFZ7tJo3A6t+2WKS6So/Q/eTcVYt2IONkpJux2ONVP2nok7wuJZ6gd1YoM9LDqLKHie0
/0EgE1kmwWpcBaBoGQsWm/D8b++bMoi8YD/F+L91OCbJ0+pboKSeaD6BhjAh4ViyukDw7rHxDX2s
SA2mcDAnPZk4F+lZD0v9mKxmXI0cn4pn5x534MpMeQnQrQSniTIrfxDkkaTXBQDk4k08rhieEep4
4pM/mx+RJPRm9dClvHSPmp+NQnv9Rt540vyiuYILbotgO9Zo/SjBgilDTAFkGBqwkMFgDQGEPUlu
rcu2vI0U6C0JvgI1m/PAB8zBgl88YAoO+bumn+b4Ua96FD4RYq95EUj0JyckMn+gHmZo4WaUtB67
VsYiOo5cqIhcCK6crmv58/ADcdnVzczaHfM4JbM+zJ5Pqn9zBKBGE8mGXjcn48lpe7vL6Mw1r+Nb
ojEf8BOh0AwVRQlRHZJSjTsurx5mMkaVxAMm6UAR+qEzOluw9jQ3Yk3U+IunOZABqFbUAuoWBtDj
AdkUxybphnVbcfWibNev3Rsmh55fQG0gMXV4y2tPEepLfPG6x4/5lhdJ5vYD5wmE19s2aUIeVDZi
OihEqyKAJP4JSH+hPEDsfG2NF/4hb6CGJ/J96kU4qpaALhU0myIGEgsPRBYdzGKp3Zxw3+5Ubhat
fxeXlTkkma9PVLaruJBpjxNraJGFKMmYnof6E99dHQRsT9VJlm9bjWI5xvgFy/V5YBFxqfH0GXzZ
qwnpXxRoC4BBqeiuolTaabNzeHerEn1Kpsxk+BH/jI0SbzIoEPF9TLf9Ky5DGrgqrK25CEmAeISq
6WUlXp6dbhxvpWUaYaDdAsKpmd+QWr+dV0t5u98ubkrzLcG3xTfjkPvVwNnMEl8h0dbJvaGJba6o
aRcCOE0qsX7ZYetESJporNKig+o+M0PCC+5UeTxHz1ZQskrX3aiaG5A+3bTU0zdWnCEwrjItMTfE
Tu6l04aSn4owdrq3aHzn5V/B8Vs5AQqTGavndET25idjlD5R1Jvs48z8FD2CpuczrPUYEkl6tNs0
TeYuwG1HsLehrwjHCPojUJgKQdmG/LWGLC1MsHDuLJlhF7pFJa3gE8VEtSV+Mu6gysv9fowUBhbr
OQ4m23N8BpLwlhq64tmIZ5kEYrGCg91Q1Q9BJ66S9eCaM5G/3I1gMplqputwS9hn6FsFB6YBBG41
6bJrW/xCByAb2ih4qQ6h9WqJVXbuDSA+cSzn83fpKterRR1f5Dt9DJJhIIXRpAOV4X/DbX038O2c
jb19Q7M9Ek7jPlvMpzY+ScF7F5MiAVA5RgayycNz0K1gCKPcYraiTv7GcdC8FTjnJFyi1Vkqe1yl
hDGVzCB/ucOPRJPoVv6knQXpFdXH+j8LA9luZUfw/4yLJ1ZgdbjHybrfmXXkjcOFiZgtrTYN9HLY
VbyKcjD5f/qIL9gKxihEm+oWRL+G7dt7z0pUAem5zsZWgpmk+EhiTvaoHgd+xKB8jANgAS74Kj/n
9OtJcZRS3XKihN/e7LtwkDRjqyeeoLVimtscH7eClRXO4pLHUeYsNZfUdCK0TGqpEr87X6UGOxMU
1czghuOn5BLBGRuOZxQtWJb9GEV/mn1zm5nrjtszix21NXgegFXH8/qgqWFAOiH++OHylkFOm7dt
TIYJM+z6W3G0DL5+ylxT3b+tdzr+J0liqfhTYHZGGVAuyslKUBgluvV4+Q+bkoYXxZqDdgfraP3y
xN6AAipvn9pOXmzIZyhiwjsfjRq8MOc6FA4d52OkK3a4AOGuDL/V/i/FA+EnSd/rXS/pOlaCBay5
PdZMl34idWBPuVa8MsueuCyVn+lzLzLbd0cUP3wt6im5sUyJ0DqqUXHABaLkLbWZY/vTjTT1yIyn
8oDxrQstboqApL7VfCgqpPTpJcSXy9CZvqxWAaH8Xp75vgPQp8z5p1OkO40PhzX9nCTbaauSY1Pv
+0AAUvl45QBXFnh8kz5IRMHjvPJi4rUtTkuq8ZIBkH6d6wsAStbFrSFlZp0lnovFSWGm466OqDdx
RHkOrlUw7I1fgtjC2xWvyqFE87aiZlFlk6CYzt3rMXFRtPFZOFMp/36lSr3c76yjnPPFm7kqw2G8
ReTAv8EUYz9ViYYr86HppuJzP88Knv4bQddwy/bPCX4ae5dO48yKJDfFSqUW443NKuuP/1k3Nds4
jqJyr1zdzNLAlVaE4ShfvUBwOI6tCY94yaImtDY6hriOernqHlm4XM2FPV2V1JG1NATQOZh815W6
HPmEAj9KGxJ/xLJjO1PA0GyBegW66GdcHrv5LalnIZZkzkNHhn9vjhsaCbKMT2q8KEHImwf1VCuV
xGaXh/EJDFbCqNS810D8F6NAekmIjp8KC+FMh9i7neZs1KP2p6pon3OALcJdrIhESliv8MeN51wI
5Zlyk9EmJ4a7BCLSxj4i2DJExf3J8vIgi24lbbWZpZE4e0FsrhbebgE8G1paRXtY10TfiSAr/UFX
9eDkCyNPO1Tz3kEIpGf7GyOrQuv8MutisCRbWkl2JZLpcTOCvlO1kTQD2KUnpdS7vZgsw4HsUOn9
SEDKtlft7hT5WqnZoez3gNs4KOAUWLMOd6ShS8kipXvlD3DidseQ3AvkZcgajElRHLvSlz1yBhfQ
Z1ShWwWbmVCB1Zh0GkKUntTjzt2nJMjX5rvV4W2bTK9OJFr4vXhKjsQviuR+cCPP5cnk3+TUCpRA
Oc0Ykqx7rcyJrnkecKVvjj58mYlVe4irZAjTA5dKloMKMbmfxHN2N2ilOMjqTd9HHPX4dXpBmbm7
I7R0K6ugi5g5aPI873C0PmVRNEncQKVsiHzQAFjcxA8aya6Fsai94Z4yHbtxTxSfxb/h5iGdHtUg
n71yaxxIAr2PBAYAykZ/uCKiDzp9zA6VrbedqaQgoXGyqXpdhMW9k4oHudPC0y763xmNcPx4w3RY
7OpalGUlidDfMqEYZ93vHKNwYWfWtZUhvlDRHS/3LZewnHjZHf9qR4L/bsKiFbt45uDylRj2IZPC
nPm7d5xLRpYaUZZU1dHD2R9xajJeGv+edlMWCnlBlQCqLq3T8NW0BIxfcUelzQTAa+91z0ht55pV
AY6YOGy7S6tuFTnirZ7Q0+U52+Za/ZiwfzbOTEejibbJcThQg8bJh5oJwq8cIZTkg6rXUqqC6MEE
N1EjqfZVgXndvfS8OtHbvW27aEh5rRmzwBJ7ItPJAKhnRCKJ+ElChL7/qcZjUMaPoPzRpHywv4eq
9vaJ19X5hQZPfWcnjeLwJeuNEFz4TNoJ0pGv9DWAhKoVtaU6OnotuYX/taaVGJ+jvpm7t4XwxrjR
jkVnYgBQz5irrL74aegGxrKnRB8q5Aj0Oxg1T/VlMBecrgEunCzm9Y60TEnP0mcKN/mjT0f+ypg6
iMFe8o98AmpVkLXn/OHFN0sGNplxLeshgBGoA4EiG1SgDo/W48HI9nOumvU2qwLYEl+NvhgjpWcH
UAUBtoNd7hQKrwkeSgL9YP1xgTHYvrQLc4uN2D3gGFDoK1M242YtGMX/33j06vqzrjtAEeSM7rni
NE7OUmmxNmpzlZl9Y0B+zOtaW3GSkWK31AEggDtMMKo+qEqq63WboLLbl6G2HyeSOgPhwZ/x1sQf
fHphNuuWqCYuo8Xv8Qgm2MDO7ijoghG7IDLfdl2L+4NbTiJMM3CszFMGrQXoE1HM/gYtW8xqRo5k
yYU1FtY01DSnlVye8E2bPy1mj04GwjK3dprZ+BiE9HbEpPsNnylDiO1ZOTzBtNa3/4eXSGBy43Hp
rE+Y3yNOtvX3w/g3Nera7yhajub9uEMf9cLI3lgAWUajQCLnk0yS/oasfvN0DYB1zbI1FB+DHqzN
3lrd87ajFt+WmkmugIppj0Q6nJuA+qi6Ok556DsRbbkOD60FQRZT7wTPJjJhzZ6ijSDzuORFy508
6x2gqPYsMCg7BAe4b6sZs+C5ducH/VNkbtuV7E6sFzGiu4a0k74E6Yxdt8o3RK/AzaUybggx21VY
akN9KWayN62BYkU42khmIAIYjbwlYn06aQ1o72Jz+gWKDaCJyaKw1s5sROIEijU6/0H7B2hYynxx
PLpM5kWEiMFgLnn5kmZsL5axm/Ys65CAGnXdfn//nrNu6+YHGhQGkQMQyr/9WlSWCXJWJ+JbshpC
BrYahYC9Ldrmh8d1lWu1Biy1OsVKb9F1cEBkbmCg7qH79HSdAvNfTC2jNK9m9SS9I2xmGrAhe1Zn
ZHrwE/6hyAaplAcwsXeMcPsM4l/oVGnWg/x/LQPG7oGDxosooGsZ5KWG98+MD8BwBpjuXPAPud29
sXqGoUrtWktcUM4jBAhCY5lStNi6akXNQ/IMhGd6NSnsuSDTCPidBt5a9WVFanAKprebb7EMU2pn
CTltqhpSjJ4H9i6YU1bZTdtgPpkrhUD6q+KZJWCGzQgkwU1KHkz4U8i8Q1Cql/GrHzurFmpOJmv9
vn562/F/eEWP9HfMKaasVC0iJX8UiYGt+iNfm4TUnXmrM1hBBbHX/Kit9JwqrJ3wFXN+zr/lE+7W
9s0/BmKcHAiqP8QB3zIpN7FCRF0AYBBZp5bwOermDXCMPZp+/81stB2Qv99VwXjT4qn3C8f9Acy0
wJyMDxYJSi/GCv5yXyUC0txW6A1IEY6m3N/J7LUtVfeIaTuDb0XhbbXUUQdRVWKX5GJKzGJngEA3
bGYgV/Kuvik1XsNn2Re4/jkC+WgGfmBNiVH2Sr5qwOhXs/+nyRG1U0WM5or0n48PYRzO0s1Otrlx
JWTK6EMHREuGlkQgLclm1ttQrf7j170mern4Qm6bf2iNzv+0Ul0uAZiz4HK2gWgou9xQ94usuGBj
qzpIwgrSTQSjqW7RhlhUQdB6g8Ycv94ZV835wxrTr2bpye466UjiIcCHD+ZRwBF51Ri6WuQpzqPx
/jxskCE5lxXnOj462QQMdcBbwkKhhIcBPYvyHgldPBWbHOGsBvWFIyz2KK/9LHlI1EsNF9kC7zyf
PtES3a04IGRhtj4HduRvK1CzTdHS0hnJcdbPrNSsfLbTXU5DjMXZNm9Fz+4ascQH7AKyPeRBwXkh
lR9bpdnU1w7BfMoqRzrq1XOGPmflUwES0QyvT6LMzt+/Kkb1WSWf+iZhIGwgjmF/Dlr3z8TDMN1L
SZoXl6Rz9311zJsWK+3Ht/ebAe5NkHIx14KSxtH7FdEn7KKpZh1zZ0SqEJxqQ+fANy9nUuG+qWPQ
Q0X/B388QryApyBFN2NvQ1BcOCiKA6sQqnKS/4W9ZFMxdGMslOg7ywE45C/HDyzsRIy+o3ui8TsW
A494CyK5mV8XSnif2P2kcXipfn0p2O2+dRlcVwGbTCphBWp/UVidGt5QHMLvz+MGcXwHxjCSws1v
Rdp1fJ231IcH0coEOnGOS0Vn+dqFAo6oXm7w0PFjFSjFtF75CjQiWzG1zbSyVZ1ZTUciO86rmMsT
e7Yih/en4jTTnX8KEw2TQGLWDwIAyEhou8GQ/NMlDplC70UuAVnfRVIZmAUFlVF5dCqP9z9D711f
jHllKFv0ansrY+aJQlyklaCEIxPya1Kc/4lWVuazZnye+U1hZzWFlRYoOJOJROQR3T7Lsi3j/bPk
SGSju74hnbPNxt30Fxa06dRF7537+vA18+TTeq26hJJT1l2LHrtkZ5z1l2ymPDIZnCmRVIRAcVZZ
CuwkZutiZF7y86Wy+2yNVNtqaDmcZlE90PCy7O5n63eHFIsK5kQFBTwAynrCWlTSjH840TCi7OCC
S87mOkMF8hBwmhJRjYhZarO9m1GNZiOaRUe6+2cx280tLIl1jcxauQV5SyToc+wgYlrJ8t6w/cGK
D1zKd8/DxQXwhK0QW4EYkckw7QFjz1IVXzAtfQjQQLipShYpJPZbLvwZ2SbB23uAFgClILVruwyK
HPSeaZBA/NcuzNQO68g4QlGgjiIM1eQbtAB+PMmQJyQw9fDd5+vTC3sIca7yPt3Kdvv37Ow2SDEp
ynsNjrl6IqGpEWEBwan1nOPGYta+VzNW4dFcxI75/hEPrHQY5wbAef3GppxuO7B6CQ8P2NtRw6dr
29pdWTuFCCQVnb1CSGi5U7mnON02WaaxR4gtZItB1Z3OkV8u0vjRHfOfGZvYDTcc2Z7fDtb+ApoR
dPMjOR09QN+0xX/AfLRa8ys/t4GZbS/UEFPp00WCx0ONM2x1KagyUyl02jRI01t96Aui/y/zUvO6
F+ZFXn20F5/XqukTCJZAEZUX10giIpD8hthAP01B4RQgMspdg4AqX1fu8uqCvelQHPclBKygn6re
eVnpqfz6Bk7cp7c+kLQOqUlgYrb+DreXRvfUweSgbtsgAaYBZkM2l3gdcilTjSk3nSDY1HI7F5Rh
MvuwfSeoX/GpNrSbcsnjMJXduVDYVIYtEvBMMhuOAsdkA0EvqDkFNkMDZ8m/6VNF+1SlqI2bWxPt
nFfK+S5jKcWjInANhFh/MElrZm3ONL6tH++6H9cKjBf+htWOGj09HjBcPBxMrvTD5A44mOCdT8Eg
6gy/hGDk5bKotBOHrVz/SNrP2sl9zEVjpSpV1a/tbkI+6ghdnYYZE2+YLmX1jY+liCohUkhWliRQ
zeLXtHhD1EK1+mHispQuyHj3oBvChrgEWniMtdCEgh6LmFtoWQk+EqE0HJeqj0zKME/6MwnmUT5X
OTS1TqqskO4u3k+atwnOCReoXpyJfXP0SpyQ8nuSCn7c0RfGEi79lsTidZU12SsABS+iKXzZq8js
v+tgFKuRyp0mF2BmolndQAnQAguMUEuHKmwVmcI3CGxFCinWMWAOdVDSxELh5o3ETwU7LwmrxMD2
fbSQNfhx5xBEpzuXSkWRiK2ffntbJLwjQY8edM2P6Z05y6kHah9Nsjg994WpszsMgSwlkXEXKRKO
iHLpZqNJjY0gYpIXWOt6xEJ/RC7niLXSYqXS0OtlsLneRrcsT94Q8JqUTqOTa/sHmw/ehMn0izuN
1KLRol7DRjtfrjMrDR3tjK8+oYkZK+NT664WfXpLub74jJjIh9GQbnoC6VI8ggY7WT80fXgqkBWp
pmc5uvLl5IYiqDVTwYnpcAE/25pQguK8xaz3NSTBCtMunpdo34iBeyNoAI1ubpvZpNas313GwWOL
4xcTNqAR0/U39q4BhoPLZGBMYGqWkHFBE4ESUjZn5/+cQjGRFPreAJaCNDKWslCJXqyRIspT1CC0
B7YLjj8Tn+gsdNPMnhAdDf/zbKspzlZ7CxciPxcdetHRdCnILCFzHRD44fnJAmBK8mtF4m4Fen/H
2Ggq5sl3hV1ziTy6De5WHQ7pPDHZJkZPIP+ljBh7z9/bLtWKFBAvWuhsErUaXKa+LvEkjQSCrS/C
L0hABqQmR1Zhh9fBoMbqNP+KfwKQ7Drja8BGbi06jmsHPIYDYqQo7V3NlSOheV7s4Z1y4pewbJlp
Ph75JJt7axbmUVbF4H3rOLDRbPd0VwdR7lBnfOFHBq2NbYWG0aiXvj4PmD5pSKpf2BeTJDFkX/AI
u34CiLx7WuthskxI1zB5Gx+zXcqLgp8rH7Ag5W1lgh1EtjdxnAvufvskeW1oQovaVghMj0bapvqL
lAPZQXw3altG1QAIS8OtgT96r+NVfXuPVJGDM165Pv01djLyoYBZaUJvxgYvycoOe/FqYCSYiUtN
D5X2CvwEtkR/vwBP+N3/0Oap3hkenJHFjF+X/mDDJLzhVAJzG5MuckMQynVtXarwLbkVJ5s3wvGI
fx2dnOIe
`pragma protect end_protected
