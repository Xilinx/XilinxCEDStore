.GT_REFCLK0(gt_refclk0_out),

.apb3clk(iffctrlq2apb3clk),
.axisclk(iffctrlq2axisclk),

.apb3psel(iffctrlq2psel),
.apb3paddr(iffctrlq2paddr),
.apb3prdata(iffctrlq2prdata),
.apb3pready(iffctrlq2pready),
.apb3pwdata(iffctrlq2pwdata),
.apb3pwrite(iffctrlq2pwrite),
.apb3penable(iffctrlq2penable),
.apb3presetn(iffctrlq2presetn),
.apb3pslverr(iffctrlq2pslverr),

.bgpdb(iffctrlq2bgpwrdnb),
.bgbypassb(iffctrlq2bgbypass),
.bgrcalovrd(iffctrlq2bgrcalctl),
.bgmonitorenb(iffctrlq2bgtesten),
.bgrcalovrdenb(iffctrlq2bgrcalovrdenb),

.ch0_rxdata(iffcq20rxdata),
.ch0_rxrate(iffcq20rxrate),
.ch0_txdata(iffcq20txdata),
.ch0_txrate(iffcq20txrate),
.ch0_bufgtce(iffcq20bufgtce),
.ch0_gtrsvd(iffcq20pinrsrvd),
.ch0_pcierstb(iffcq20perstb),
.ch0_rxctrl0(iffcq20rxctrl0),
.ch0_rxctrl1(iffcq20rxctrl1),
.ch0_rxctrl2(iffcq20rxctrl2),
.ch0_rxctrl3(iffcq20rxctrl3),
.ch0_rxlpmen(iffcq20rxlpmen),
.ch0_rxpkdet(q2_ch0_rxpkdet),
.ch0_rxqpien(iffcq20rxqpien),
.ch0_rxslide(iffcq20rxslide),
.ch0_rxvalid(iffcq20rxvalid),
.ch0_tstclk0(iffcq20tstclk0),
.ch0_tstclk1(iffcq20tstclk1),
.ch0_txctrl0(iffcq20txctrl0),
.ch0_txctrl1(iffcq20txctrl1),
.ch0_txctrl2(iffcq20txctrl2),
.ch0_txpippmen(iffcq20enppm),
.ch0_txswing(iffcq20txswing),
.ch0_rxpd(iffcq20rxpowerdown),
.ch0_txpd(iffcq20txpowerdown),
.ch0_bufgtdiv(iffcq20bufgtdiv),
.ch0_bufgtrst(iffcq20bufgtrst),
.ch0_iloreset(iffcq20iloreset),
.ch0_loopback(iffcq20loopback),
.ch0_phyready(iffcq20phyready),
.ch0_rxcdrhold(iffcq20cdrhold),
.ch0_rxcdrlock(iffcq20cdrlock),
.ch0_rxheader(iffcq20rxheader),
.ch0_rxlatclk(iffcq20rxlatclk),
.ch0_rxoutclk(q2_ch0_rxoutclk),
.ch0_rxstatus(iffcq20rxstatus),
.ch0_rxusrclk(iffcq20rxusrclk),
.ch0_txcomsas(iffcq20txcomsas),
.ch0_txdeemph(iffcq20txdeemph),
.ch0_txheader(iffcq20txheader),
.ch0_txlatclk(iffcq20txlatclk),
.ch0_txmargin(iffcq20txmargin),
.ch0_txoutclk(q2_ch0_txoutclk),
.ch0_txusrclk(iffcq20txusrclk),
.ch0_dfehold(iffcq20aptexthold),
.ch0_rxuserrdy(iffcq20rxusrrdy),
.ch0_txuserrdy(iffcq20txusrrdy),
.ch0_cdrfreqos(iffcq20cdrfreqos),
.ch0_cdrstepsq(iffcq20cdrstepsq),
.ch0_cdrstepsx(iffcq20cdrstepsx),
.ch0_dfeovrd(iffcq20aptoverwren),
.ch0_dmonitorclk(iffcq20dmonclk),
.ch0_dmonitorout(iffcq20dmonout),
.ch0_gtrxreset(iffcq20gtrxreset),
.ch0_gttxreset(iffcq20gttxreset),
.ch0_pcsrsvdin(iffcq20pcsrsvdin),
.ch0_phystatus(iffcq20phystatus),
.ch0_rxchbondi(iffcq20rxchbondi),
.ch0_rxchbondo(iffcq20rxchbondo),
.ch0_rxprbserr(iffcq20rxprbserr),
.ch0_rxprbssel(iffcq20rxprbssel),
.ch0_rxqpisenn(iffcq20rxqpisenn),
.ch0_rxqpisenp(iffcq20rxqpisenp),
.ch0_txcominit(iffcq20txcominit),
.ch0_txcomwake(iffcq20txcomwake),
.ch0_txdccdone(iffcq20txdccdone),
.ch0_txdiffctrl(iffcq20txdrvamp),
.ch0_txinhibit(iffcq20txinhibit),
.ch0_txpisopd(iffcq20txserpwrdn),
.ch0_txprbssel(iffcq20txprbssel),
.ch0_txqpisenn(iffcq20txqpisenn),
.ch0_txqpisenp(iffcq20txqpisenp),
.ch0_clkrsvd0(iffcq20ckpinrsrvd0),
.ch0_clkrsvd1(iffcq20ckpinrsrvd1),
.ch0_pinrsvdas(iffcq20pinrsrvdas),
.ch0_rxcdrovrden(iffcq20cdrovren),
.ch0_rxosintdone(iffcq20cfokdone),
.ch0_txprecursor(iffcq20txemppre),
.ch0_cdrstepdir(iffcq20cdrstepdir),
.ch0_pcsrsvdout(iffcq20pcsrsvdout),
.ch0_refdebugout(iffcq20refclkpma),
.ch0_rxcdrreset(iffcq20cdrphreset),
.ch0_rxcommadet(iffcq20rxcommadet),
.ch0_rxcomsasdet(iffcq20comsasdet),
.ch0_rxelecidle(iffcq20rxelecidle),
.ch0_rxoobreset(iffcq20rxoobreset),
.ch0_rxpolarity(iffcq20rxpolarity),
.ch0_rxsliderdy(iffcq20rxsliderdy),
.ch0_rxslipdone(iffcq20rxslipdone),
.ch0_rxsyncdone(iffcq20rxsyncdone),
.ch0_txelecidle(iffcq20txelecidle),
.ch0_txpolarity(iffcq20txpolarity),
.ch0_txpostcursor(iffcq20txemppos),
.ch0_txsequence(iffcq20txsequence),
.ch0_txsyncdone(iffcq20txsyncdone),
.ch0_cdrbmcdrreq(iffcq20cdrbmcdreq),
.ch0_rxclkcorcnt(iffcq20rxckcorcnt),
.ch0_txmaincursor(iffcq20txempmain),
.ch0_bufgtcemask(iffcq20bufgtcemask),
.ch0_cdrincpctrl(iffcq20cdrincpctrl),
.ch0_rxbufstatus(iffcq20rxbufstatus),
.ch0_rxcdrphdone(iffcq20rxcdrphdone),
.ch0_rxcominitdet(iffcq20cominitdet),
.ch0_rxcomwakedet(iffcq20comwakedet),
.ch0_rxdapireset(iffcq20rxdapireset),
.ch0_rxdatavalid(iffcq20rxdatavalid),
.ch0_rxresetdone(iffcq20rxresetdone),
.ch0_rxresetmode(iffcq20rxresetmode),
.ch0_rxsyncallin(iffcq20rxsyncallin),
.ch0_txbufstatus(iffcq20txbufstatus),
.ch0_txcomfinish(iffcq20txcomfinish),
.ch0_txdapireset(iffcq20txdapireset),
.ch0_txoneszeros(iffcq20txoneszeros),
.ch0_txqpibiasen(iffcq20txqpibiasen),
.ch0_txqpiweakpu(iffcq20txqpiweakpu),
.ch0_txresetdone(iffcq20txresetdone),
.ch0_txresetmode(iffcq20txresetmode),
.ch0_txsyncallin(iffcq20txsyncallin),
.ch0_rxphdlypd(iffcq20rxphasealignpd),
.ch0_txphdlypd(iffcq20txphasealignpd),
.ch0_bufgtrstmask(iffcq20bufgtrstmask),
.ch0_eyescanreset(iffcq20eyescanreset),
.ch0_hsdppcsreset(iffcq20hsdppcsreset),
.ch0_iloresetdone(iffcq20iloresetdone),
.ch0_iloresetmask(iffcq20iloresetmask),
.ch0_rxdebugpcsout(iffcq20rxoutpcsclk),
.ch0_rxeqtraining(iffcq20rxeqtraining),
.ch0_rxphdlyreset(iffcq20rxphdlyreset),
.ch0_rxprbslocked(iffcq20rxprbslocked),
.ch0_rxstartofseq(iffcq20rxstartofseq),
.ch0_txdebugpcsout(iffcq20txoutpcsclk),
.ch0_txphdlyreset(iffcq20txphdlyreset),
.ch0_rxmstreset(iffctrlq2mstrxreset[0]),
.ch0_txmstreset(iffctrlq2msttxreset[0]),
.ch0_dmonfiforeset(iffcq20dmonfiforeset),
.ch0_rx10gstat(iffcq20rxethernetstatout),
.ch0_rxbyterealign(q2_ch0_rxbyterealign),
.ch0_rxchanbondseq(iffcq20rxchanbondseq),
.ch0_rxchanrealign(iffcq20rxchanrealign),
.ch0_rxgearboxslip(iffcq20rxgearboxslip),
.ch0_rxheadervalid(iffcq20rxheadervalid),
.ch0_rxmldchainreq(iffcq20rxmldchainreq),
.ch0_rxtermination(iffcq20rxtermination),
.ch0_txmldchainreq(iffcq20txmldchainreq),
.ch0_txpippmstepsize(iffcq20stepsizeppm),
.ch0_txswingoutlow(iffcq20txswingoutlow),
.ch0_rxphalignerr(iffcq20rxphasealignerr),
.ch0_rxphalignreq(iffcq20rxphasealignreq),
.ch0_txphalignerr(iffcq20txphasealignerr),
.ch0_txphalignreq(iffcq20txphasealignreq),
.ch0_txphdlytstclk(iffcq20tcoclkfsmfrout),
.ch0_dmonitoroutclk(q2_ch0_dmonitoroutclk),
.ch0_eyescantrigger(iffcq20eyescantrigger),
.ch0_resetexception(iffcq20resetexception),
.ch0_rxchanisaligned(iffcq20rxchisaligned),
.ch0_rxdlyalignerr(iffcq20rxdelayalignerr),
.ch0_rxdlyalignreq(iffcq20rxdelayalignreq),
.ch0_rxmldchaindone(iffcq20rxmldchaindone),
.ch0_rxpcsresetmask(iffcq20rxpcsresetmask),
.ch0_rxpmaresetdone(iffcq20rxpmaresetdone),
.ch0_rxpmaresetmask(iffcq20rxpmaresetmask),
.ch0_rxprbscntreset(iffcq20rxprbscntreset),
.ch0_rxprogdivreset(iffcq20rxprogdivreset),
.ch0_txdetectrx(iffcq20txdetectrxloopback),
.ch0_txdlyalignerr(iffcq20txdelayalignerr),
.ch0_txdlyalignreq(iffcq20txdelayalignreq),
.ch0_txmldchaindone(iffcq20txmldchaindone),
.ch0_txpcsresetmask(iffcq20txpcsresetmask),
.ch0_txpicodereset(iffcq20txtxpicodereset),
.ch0_txpmaresetdone(iffcq20txpmaresetdone),
.ch0_txpmaresetmask(iffcq20txpmaresetmask),
.ch0_txprbsforceerr(iffcq20txprbsforceerr),
.ch0_txprogdivreset(iffcq20txprogdivreset),
.ch0_txswingouthigh(iffcq20txswingouthigh),
.ch0_rxphaligndone(iffcq20rxphasealigndone),
.ch0_txphaligndone(iffcq20txphasealigndone),
.ch0_rxbyteisaligned(iffcq20rxbyteisaligned),
.ch0_rxdapicodereset(iffcq20rxdapicodereset),
.ch0_rxdapiresetdone(iffcq20rxdapiresetdone),
.ch0_rxdapiresetmask(iffcq20rxdapiresetmask),
.ch0_rxfinealigndone(iffcq20rxfinealigndone),
.ch0_rxphshift180(iffcq20rxphaseshift180req),
.ch0_txdapicodereset(iffcq20txdapicodereset),
.ch0_txdapiresetdone(iffcq20txdapiresetdone),
.ch0_txdapiresetmask(iffcq20txdapiresetmask),
.ch0_txphalignoutrsvd(iffcq20txchicooutrsvd),
.ch0_txphshift180(iffcq20txphaseshift180req),
.ch0_txpicodeovrden(iffcq20txtxpicodeovrden),
.ch0_rxphsetinitreq(iffcq20rxphasesetinitreq),
.ch0_txphsetinitreq(iffcq20txphasesetinitreq),
.ch0_eyescandataerror(iffcq20eyescandataerror),
.ch0_rxdapicodeovrden(iffcq20rxdapicodeovrden),
.ch0_rxmlfinealignreq(iffcq20rxmlfinealignreq),
.ch0_txdapicodeovrden(iffcq20txdapicodeovrden),
.ch0_rxmstresetdone(iffctrlq2mstrxresetdone[0]),
.ch0_rxphsetinitdone(iffcq20rxphasesetinitdone),
.ch0_txmstresetdone(iffctrlq2msttxresetdone[0]),
.ch0_txphsetinitdone(iffcq20txphasesetinitdone),
.ch0_rxdlyalignprog(iffcq20rxdelayalignprogress),
.ch0_rxphalignresetmask(iffcq20rxchicoresetmask),
.ch0_txdlyalignprog(iffcq20txdelayalignprogress),
.ch0_txpausedelayalign(iffcq20txpausedelayalign),
.ch0_txphalignresetmask(iffcq20txchicoresetmask),
.ch0_xpipe5_pipeline_en(iffcq20xpipe5pipelineen),
.ch0_phyesmadaptsave(iffcq20phyesmadaptationsave),
.ch0_rxphshift180done(iffcq20rxphaseshift180done),
.ch0_tx10gstat(iffcq20txethernetstattxlocalfault),
.ch0_txphshift180done(iffcq20txphaseshift180done),
.ch0_rxprogdivresetdone(iffcq20rxprogdivresetdone),
.ch0_rxsimplexphystatus(iffcq20rxsimplexphystatus),
.ch0_txprogdivresetdone(iffcq20txprogdivresetdone),
.ch0_txsimplexphystatus(iffcq20txsimplexphystatus),
.ch0_rxphdlyresetdone(iffcq20rxphasedelayresetdone),
.ch0_txphdlyresetdone(iffcq20txphasedelayresetdone),

.ch1_rxdata(iffcq21rxdata),
.ch1_rxrate(iffcq21rxrate),
.ch1_txdata(iffcq21txdata),
.ch1_txrate(iffcq21txrate),
.ch1_bufgtce(iffcq21bufgtce),
.ch1_gtrsvd(iffcq21pinrsrvd),
.ch1_pcierstb(iffcq21perstb),
.ch1_rxctrl0(iffcq21rxctrl0),
.ch1_rxctrl1(iffcq21rxctrl1),
.ch1_rxctrl2(iffcq21rxctrl2),
.ch1_rxctrl3(iffcq21rxctrl3),
.ch1_rxlpmen(iffcq21rxlpmen),
.ch1_rxpkdet(q2_ch1_rxpkdet),
.ch1_rxqpien(iffcq21rxqpien),
.ch1_rxslide(iffcq21rxslide),
.ch1_rxvalid(iffcq21rxvalid),
.ch1_tstclk0(iffcq21tstclk0),
.ch1_tstclk1(iffcq21tstclk1),
.ch1_txctrl0(iffcq21txctrl0),
.ch1_txctrl1(iffcq21txctrl1),
.ch1_txctrl2(iffcq21txctrl2),
.ch1_txpippmen(iffcq21enppm),
.ch1_txswing(iffcq21txswing),
.ch1_rxpd(iffcq21rxpowerdown),
.ch1_txpd(iffcq21txpowerdown),
.ch1_bufgtdiv(iffcq21bufgtdiv),
.ch1_bufgtrst(iffcq21bufgtrst),
.ch1_iloreset(iffcq21iloreset),
.ch1_loopback(iffcq21loopback),
.ch1_phyready(iffcq21phyready),
.ch1_rxcdrhold(iffcq21cdrhold),
.ch1_rxcdrlock(iffcq21cdrlock),
.ch1_rxheader(iffcq21rxheader),
.ch1_rxlatclk(iffcq21rxlatclk),
.ch1_rxoutclk(q2_ch1_rxoutclk),
.ch1_rxstatus(iffcq21rxstatus),
.ch1_rxusrclk(iffcq21rxusrclk),
.ch1_txcomsas(iffcq21txcomsas),
.ch1_txdeemph(iffcq21txdeemph),
.ch1_txheader(iffcq21txheader),
.ch1_txlatclk(iffcq21txlatclk),
.ch1_txmargin(iffcq21txmargin),
.ch1_txoutclk(q2_ch1_txoutclk),
.ch1_txusrclk(iffcq21txusrclk),
.ch1_dfehold(iffcq21aptexthold),
.ch1_rxuserrdy(iffcq21rxusrrdy),
.ch1_txuserrdy(iffcq21txusrrdy),
.ch1_cdrfreqos(iffcq21cdrfreqos),
.ch1_cdrstepsq(iffcq21cdrstepsq),
.ch1_cdrstepsx(iffcq21cdrstepsx),
.ch1_dfeovrd(iffcq21aptoverwren),
.ch1_dmonitorclk(iffcq21dmonclk),
.ch1_dmonitorout(iffcq21dmonout),
.ch1_gtrxreset(iffcq21gtrxreset),
.ch1_gttxreset(iffcq21gttxreset),
.ch1_pcsrsvdin(iffcq21pcsrsvdin),
.ch1_phystatus(iffcq21phystatus),
.ch1_rxchbondi(iffcq21rxchbondi),
.ch1_rxchbondo(iffcq21rxchbondo),
.ch1_rxprbserr(iffcq21rxprbserr),
.ch1_rxprbssel(iffcq21rxprbssel),
.ch1_rxqpisenn(iffcq21rxqpisenn),
.ch1_rxqpisenp(iffcq21rxqpisenp),
.ch1_txcominit(iffcq21txcominit),
.ch1_txcomwake(iffcq21txcomwake),
.ch1_txdccdone(iffcq21txdccdone),
.ch1_txdiffctrl(iffcq21txdrvamp),
.ch1_txinhibit(iffcq21txinhibit),
.ch1_txpisopd(iffcq21txserpwrdn),
.ch1_txprbssel(iffcq21txprbssel),
.ch1_txqpisenn(iffcq21txqpisenn),
.ch1_txqpisenp(iffcq21txqpisenp),
.ch1_clkrsvd0(iffcq21ckpinrsrvd0),
.ch1_clkrsvd1(iffcq21ckpinrsrvd1),
.ch1_pinrsvdas(iffcq21pinrsrvdas),
.ch1_rxcdrovrden(iffcq21cdrovren),
.ch1_rxosintdone(iffcq21cfokdone),
.ch1_txprecursor(iffcq21txemppre),
.ch1_cdrstepdir(iffcq21cdrstepdir),
.ch1_pcsrsvdout(iffcq21pcsrsvdout),
.ch1_refdebugout(iffcq21refclkpma),
.ch1_rxcdrreset(iffcq21cdrphreset),
.ch1_rxcommadet(iffcq21rxcommadet),
.ch1_rxcomsasdet(iffcq21comsasdet),
.ch1_rxelecidle(iffcq21rxelecidle),
.ch1_rxoobreset(iffcq21rxoobreset),
.ch1_rxpolarity(iffcq21rxpolarity),
.ch1_rxsliderdy(iffcq21rxsliderdy),
.ch1_rxslipdone(iffcq21rxslipdone),
.ch1_rxsyncdone(iffcq21rxsyncdone),
.ch1_txelecidle(iffcq21txelecidle),
.ch1_txpolarity(iffcq21txpolarity),
.ch1_txpostcursor(iffcq21txemppos),
.ch1_txsequence(iffcq21txsequence),
.ch1_txsyncdone(iffcq21txsyncdone),
.ch1_cdrbmcdrreq(iffcq21cdrbmcdreq),
.ch1_rxclkcorcnt(iffcq21rxckcorcnt),
.ch1_txmaincursor(iffcq21txempmain),
.ch1_bufgtcemask(iffcq21bufgtcemask),
.ch1_cdrincpctrl(iffcq21cdrincpctrl),
.ch1_rxbufstatus(iffcq21rxbufstatus),
.ch1_rxcdrphdone(iffcq21rxcdrphdone),
.ch1_rxcominitdet(iffcq21cominitdet),
.ch1_rxcomwakedet(iffcq21comwakedet),
.ch1_rxdapireset(iffcq21rxdapireset),
.ch1_rxdatavalid(iffcq21rxdatavalid),
.ch1_rxresetdone(iffcq21rxresetdone),
.ch1_rxresetmode(iffcq21rxresetmode),
.ch1_rxsyncallin(iffcq21rxsyncallin),
.ch1_txbufstatus(iffcq21txbufstatus),
.ch1_txcomfinish(iffcq21txcomfinish),
.ch1_txdapireset(iffcq21txdapireset),
.ch1_txoneszeros(iffcq21txoneszeros),
.ch1_txqpibiasen(iffcq21txqpibiasen),
.ch1_txqpiweakpu(iffcq21txqpiweakpu),
.ch1_txresetdone(iffcq21txresetdone),
.ch1_txresetmode(iffcq21txresetmode),
.ch1_txsyncallin(iffcq21txsyncallin),
.ch1_rxphdlypd(iffcq21rxphasealignpd),
.ch1_txphdlypd(iffcq21txphasealignpd),
.ch1_bufgtrstmask(iffcq21bufgtrstmask),
.ch1_eyescanreset(iffcq21eyescanreset),
.ch1_hsdppcsreset(iffcq21hsdppcsreset),
.ch1_iloresetdone(iffcq21iloresetdone),
.ch1_iloresetmask(iffcq21iloresetmask),
.ch1_rxdebugpcsout(iffcq21rxoutpcsclk),
.ch1_rxeqtraining(iffcq21rxeqtraining),
.ch1_rxphdlyreset(iffcq21rxphdlyreset),
.ch1_rxprbslocked(iffcq21rxprbslocked),
.ch1_rxstartofseq(iffcq21rxstartofseq),
.ch1_txdebugpcsout(iffcq21txoutpcsclk),
.ch1_txphdlyreset(iffcq21txphdlyreset),
.ch1_rxmstreset(iffctrlq2mstrxreset[1]),
.ch1_txmstreset(iffctrlq2msttxreset[1]),
.ch1_dmonfiforeset(iffcq21dmonfiforeset),
.ch1_rx10gstat(iffcq21rxethernetstatout),
.ch1_rxbyterealign(q2_ch1_rxbyterealign),
.ch1_rxchanbondseq(iffcq21rxchanbondseq),
.ch1_rxchanrealign(iffcq21rxchanrealign),
.ch1_rxgearboxslip(iffcq21rxgearboxslip),
.ch1_rxheadervalid(iffcq21rxheadervalid),
.ch1_rxmldchainreq(iffcq21rxmldchainreq),
.ch1_rxtermination(iffcq21rxtermination),
.ch1_txmldchainreq(iffcq21txmldchainreq),
.ch1_txpippmstepsize(iffcq21stepsizeppm),
.ch1_txswingoutlow(iffcq21txswingoutlow),
.ch1_rxphalignerr(iffcq21rxphasealignerr),
.ch1_rxphalignreq(iffcq21rxphasealignreq),
.ch1_txphalignerr(iffcq21txphasealignerr),
.ch1_txphalignreq(iffcq21txphasealignreq),
.ch1_txphdlytstclk(iffcq21tcoclkfsmfrout),
.ch1_dmonitoroutclk(q2_ch1_dmonitoroutclk),
.ch1_eyescantrigger(iffcq21eyescantrigger),
.ch1_resetexception(iffcq21resetexception),
.ch1_rxchanisaligned(iffcq21rxchisaligned),
.ch1_rxdlyalignerr(iffcq21rxdelayalignerr),
.ch1_rxdlyalignreq(iffcq21rxdelayalignreq),
.ch1_rxmldchaindone(iffcq21rxmldchaindone),
.ch1_rxpcsresetmask(iffcq21rxpcsresetmask),
.ch1_rxpmaresetdone(iffcq21rxpmaresetdone),
.ch1_rxpmaresetmask(iffcq21rxpmaresetmask),
.ch1_rxprbscntreset(iffcq21rxprbscntreset),
.ch1_rxprogdivreset(iffcq21rxprogdivreset),
.ch1_txdetectrx(iffcq21txdetectrxloopback),
.ch1_txdlyalignerr(iffcq21txdelayalignerr),
.ch1_txdlyalignreq(iffcq21txdelayalignreq),
.ch1_txmldchaindone(iffcq21txmldchaindone),
.ch1_txpcsresetmask(iffcq21txpcsresetmask),
.ch1_txpicodereset(iffcq21txtxpicodereset),
.ch1_txpmaresetdone(iffcq21txpmaresetdone),
.ch1_txpmaresetmask(iffcq21txpmaresetmask),
.ch1_txprbsforceerr(iffcq21txprbsforceerr),
.ch1_txprogdivreset(iffcq21txprogdivreset),
.ch1_txswingouthigh(iffcq21txswingouthigh),
.ch1_rxphaligndone(iffcq21rxphasealigndone),
.ch1_txphaligndone(iffcq21txphasealigndone),
.ch1_rxbyteisaligned(iffcq21rxbyteisaligned),
.ch1_rxdapicodereset(iffcq21rxdapicodereset),
.ch1_rxdapiresetdone(iffcq21rxdapiresetdone),
.ch1_rxdapiresetmask(iffcq21rxdapiresetmask),
.ch1_rxfinealigndone(iffcq21rxfinealigndone),
.ch1_rxphshift180(iffcq21rxphaseshift180req),
.ch1_txdapicodereset(iffcq21txdapicodereset),
.ch1_txdapiresetdone(iffcq21txdapiresetdone),
.ch1_txdapiresetmask(iffcq21txdapiresetmask),
.ch1_txphalignoutrsvd(iffcq21txchicooutrsvd),
.ch1_txphshift180(iffcq21txphaseshift180req),
.ch1_txpicodeovrden(iffcq21txtxpicodeovrden),
.ch1_rxphsetinitreq(iffcq21rxphasesetinitreq),
.ch1_txphsetinitreq(iffcq21txphasesetinitreq),
.ch1_eyescandataerror(iffcq21eyescandataerror),
.ch1_rxdapicodeovrden(iffcq21rxdapicodeovrden),
.ch1_rxmlfinealignreq(iffcq21rxmlfinealignreq),
.ch1_txdapicodeovrden(iffcq21txdapicodeovrden),
.ch1_rxmstresetdone(iffctrlq2mstrxresetdone[1]),
.ch1_rxphsetinitdone(iffcq21rxphasesetinitdone),
.ch1_txmstresetdone(iffctrlq2msttxresetdone[1]),
.ch1_txphsetinitdone(iffcq21txphasesetinitdone),
.ch1_rxdlyalignprog(iffcq21rxdelayalignprogress),
.ch1_rxphalignresetmask(iffcq21rxchicoresetmask),
.ch1_txdlyalignprog(iffcq21txdelayalignprogress),
.ch1_txpausedelayalign(iffcq21txpausedelayalign),
.ch1_txphalignresetmask(iffcq21txchicoresetmask),
.ch1_xpipe5_pipeline_en(iffcq21xpipe5pipelineen),
.ch1_phyesmadaptsave(iffcq21phyesmadaptationsave),
.ch1_rxphshift180done(iffcq21rxphaseshift180done),
.ch1_tx10gstat(iffcq21txethernetstattxlocalfault),
.ch1_txphshift180done(iffcq21txphaseshift180done),
.ch1_rxprogdivresetdone(iffcq21rxprogdivresetdone),
.ch1_rxsimplexphystatus(iffcq21rxsimplexphystatus),
.ch1_txprogdivresetdone(iffcq21txprogdivresetdone),
.ch1_txsimplexphystatus(iffcq21txsimplexphystatus),
.ch1_rxphdlyresetdone(iffcq21rxphasedelayresetdone),
.ch1_txphdlyresetdone(iffcq21txphasedelayresetdone),

.ch2_rxdata(iffcq22rxdata),
.ch2_rxrate(iffcq22rxrate),
.ch2_txdata(iffcq22txdata),
.ch2_txrate(iffcq22txrate),
.ch2_bufgtce(iffcq22bufgtce),
.ch2_gtrsvd(iffcq22pinrsrvd),
.ch2_pcierstb(iffcq22perstb),
.ch2_rxctrl0(iffcq22rxctrl0),
.ch2_rxctrl1(iffcq22rxctrl1),
.ch2_rxctrl2(iffcq22rxctrl2),
.ch2_rxctrl3(iffcq22rxctrl3),
.ch2_rxlpmen(iffcq22rxlpmen),
.ch2_rxpkdet(q2_ch2_rxpkdet),
.ch2_rxqpien(iffcq22rxqpien),
.ch2_rxslide(iffcq22rxslide),
.ch2_rxvalid(iffcq22rxvalid),
.ch2_tstclk0(iffcq22tstclk0),
.ch2_tstclk1(iffcq22tstclk1),
.ch2_txctrl0(iffcq22txctrl0),
.ch2_txctrl1(iffcq22txctrl1),
.ch2_txctrl2(iffcq22txctrl2),
.ch2_txpippmen(iffcq22enppm),
.ch2_txswing(iffcq22txswing),
.ch2_rxpd(iffcq22rxpowerdown),
.ch2_txpd(iffcq22txpowerdown),
.ch2_bufgtdiv(iffcq22bufgtdiv),
.ch2_bufgtrst(iffcq22bufgtrst),
.ch2_iloreset(iffcq22iloreset),
.ch2_loopback(iffcq22loopback),
.ch2_phyready(iffcq22phyready),
.ch2_rxcdrhold(iffcq22cdrhold),
.ch2_rxcdrlock(iffcq22cdrlock),
.ch2_rxheader(iffcq22rxheader),
.ch2_rxlatclk(iffcq22rxlatclk),
.ch2_rxoutclk(q2_ch2_rxoutclk),
.ch2_rxstatus(iffcq22rxstatus),
.ch2_rxusrclk(iffcq22rxusrclk),
.ch2_txcomsas(iffcq22txcomsas),
.ch2_txdeemph(iffcq22txdeemph),
.ch2_txheader(iffcq22txheader),
.ch2_txlatclk(iffcq22txlatclk),
.ch2_txmargin(iffcq22txmargin),
.ch2_txoutclk(q2_ch2_txoutclk),
.ch2_txusrclk(iffcq22txusrclk),
.ch2_dfehold(iffcq22aptexthold),
.ch2_rxuserrdy(iffcq22rxusrrdy),
.ch2_txuserrdy(iffcq22txusrrdy),
.ch2_cdrfreqos(iffcq22cdrfreqos),
.ch2_cdrstepsq(iffcq22cdrstepsq),
.ch2_cdrstepsx(iffcq22cdrstepsx),
.ch2_dfeovrd(iffcq22aptoverwren),
.ch2_dmonitorclk(iffcq22dmonclk),
.ch2_dmonitorout(iffcq22dmonout),
.ch2_gtrxreset(iffcq22gtrxreset),
.ch2_gttxreset(iffcq22gttxreset),
.ch2_pcsrsvdin(iffcq22pcsrsvdin),
.ch2_phystatus(iffcq22phystatus),
.ch2_rxchbondi(iffcq22rxchbondi),
.ch2_rxchbondo(iffcq22rxchbondo),
.ch2_rxprbserr(iffcq22rxprbserr),
.ch2_rxprbssel(iffcq22rxprbssel),
.ch2_rxqpisenn(iffcq22rxqpisenn),
.ch2_rxqpisenp(iffcq22rxqpisenp),
.ch2_txcominit(iffcq22txcominit),
.ch2_txcomwake(iffcq22txcomwake),
.ch2_txdccdone(iffcq22txdccdone),
.ch2_txdiffctrl(iffcq22txdrvamp),
.ch2_txinhibit(iffcq22txinhibit),
.ch2_txpisopd(iffcq22txserpwrdn),
.ch2_txprbssel(iffcq22txprbssel),
.ch2_txqpisenn(iffcq22txqpisenn),
.ch2_txqpisenp(iffcq22txqpisenp),
.ch2_clkrsvd0(iffcq22ckpinrsrvd0),
.ch2_clkrsvd1(iffcq22ckpinrsrvd1),
.ch2_pinrsvdas(iffcq22pinrsrvdas),
.ch2_rxcdrovrden(iffcq22cdrovren),
.ch2_rxosintdone(iffcq22cfokdone),
.ch2_txprecursor(iffcq22txemppre),
.ch2_cdrstepdir(iffcq22cdrstepdir),
.ch2_pcsrsvdout(iffcq22pcsrsvdout),
.ch2_refdebugout(iffcq22refclkpma),
.ch2_rxcdrreset(iffcq22cdrphreset),
.ch2_rxcommadet(iffcq22rxcommadet),
.ch2_rxcomsasdet(iffcq22comsasdet),
.ch2_rxelecidle(iffcq22rxelecidle),
.ch2_rxoobreset(iffcq22rxoobreset),
.ch2_rxpolarity(iffcq22rxpolarity),
.ch2_rxsliderdy(iffcq22rxsliderdy),
.ch2_rxslipdone(iffcq22rxslipdone),
.ch2_rxsyncdone(iffcq22rxsyncdone),
.ch2_txelecidle(iffcq22txelecidle),
.ch2_txpolarity(iffcq22txpolarity),
.ch2_txpostcursor(iffcq22txemppos),
.ch2_txsequence(iffcq22txsequence),
.ch2_txsyncdone(iffcq22txsyncdone),
.ch2_cdrbmcdrreq(iffcq22cdrbmcdreq),
.ch2_rxclkcorcnt(iffcq22rxckcorcnt),
.ch2_txmaincursor(iffcq22txempmain),
.ch2_bufgtcemask(iffcq22bufgtcemask),
.ch2_cdrincpctrl(iffcq22cdrincpctrl),
.ch2_rxbufstatus(iffcq22rxbufstatus),
.ch2_rxcdrphdone(iffcq22rxcdrphdone),
.ch2_rxcominitdet(iffcq22cominitdet),
.ch2_rxcomwakedet(iffcq22comwakedet),
.ch2_rxdapireset(iffcq22rxdapireset),
.ch2_rxdatavalid(iffcq22rxdatavalid),
.ch2_rxresetdone(iffcq22rxresetdone),
.ch2_rxresetmode(iffcq22rxresetmode),
.ch2_rxsyncallin(iffcq22rxsyncallin),
.ch2_txbufstatus(iffcq22txbufstatus),
.ch2_txcomfinish(iffcq22txcomfinish),
.ch2_txdapireset(iffcq22txdapireset),
.ch2_txoneszeros(iffcq22txoneszeros),
.ch2_txqpibiasen(iffcq22txqpibiasen),
.ch2_txqpiweakpu(iffcq22txqpiweakpu),
.ch2_txresetdone(iffcq22txresetdone),
.ch2_txresetmode(iffcq22txresetmode),
.ch2_txsyncallin(iffcq22txsyncallin),
.ch2_rxphdlypd(iffcq22rxphasealignpd),
.ch2_txphdlypd(iffcq22txphasealignpd),
.ch2_bufgtrstmask(iffcq22bufgtrstmask),
.ch2_eyescanreset(iffcq22eyescanreset),
.ch2_hsdppcsreset(iffcq22hsdppcsreset),
.ch2_iloresetdone(iffcq22iloresetdone),
.ch2_iloresetmask(iffcq22iloresetmask),
.ch2_rxdebugpcsout(iffcq22rxoutpcsclk),
.ch2_rxeqtraining(iffcq22rxeqtraining),
.ch2_rxphdlyreset(iffcq22rxphdlyreset),
.ch2_rxprbslocked(iffcq22rxprbslocked),
.ch2_rxstartofseq(iffcq22rxstartofseq),
.ch2_txdebugpcsout(iffcq22txoutpcsclk),
.ch2_txphdlyreset(iffcq22txphdlyreset),
.ch2_rxmstreset(iffctrlq2mstrxreset[2]),
.ch2_txmstreset(iffctrlq2msttxreset[2]),
.ch2_dmonfiforeset(iffcq22dmonfiforeset),
.ch2_rx10gstat(iffcq22rxethernetstatout),
.ch2_rxbyterealign(q2_ch2_rxbyterealign),
.ch2_rxchanbondseq(iffcq22rxchanbondseq),
.ch2_rxchanrealign(iffcq22rxchanrealign),
.ch2_rxgearboxslip(iffcq22rxgearboxslip),
.ch2_rxheadervalid(iffcq22rxheadervalid),
.ch2_rxmldchainreq(iffcq22rxmldchainreq),
.ch2_rxtermination(iffcq22rxtermination),
.ch2_txmldchainreq(iffcq22txmldchainreq),
.ch2_txpippmstepsize(iffcq22stepsizeppm),
.ch2_txswingoutlow(iffcq22txswingoutlow),
.ch2_rxphalignerr(iffcq22rxphasealignerr),
.ch2_rxphalignreq(iffcq22rxphasealignreq),
.ch2_txphalignerr(iffcq22txphasealignerr),
.ch2_txphalignreq(iffcq22txphasealignreq),
.ch2_txphdlytstclk(iffcq22tcoclkfsmfrout),
.ch2_dmonitoroutclk(q2_ch2_dmonitoroutclk),
.ch2_eyescantrigger(iffcq22eyescantrigger),
.ch2_resetexception(iffcq22resetexception),
.ch2_rxchanisaligned(iffcq22rxchisaligned),
.ch2_rxdlyalignerr(iffcq22rxdelayalignerr),
.ch2_rxdlyalignreq(iffcq22rxdelayalignreq),
.ch2_rxmldchaindone(iffcq22rxmldchaindone),
.ch2_rxpcsresetmask(iffcq22rxpcsresetmask),
.ch2_rxpmaresetdone(iffcq22rxpmaresetdone),
.ch2_rxpmaresetmask(iffcq22rxpmaresetmask),
.ch2_rxprbscntreset(iffcq22rxprbscntreset),
.ch2_rxprogdivreset(iffcq22rxprogdivreset),
.ch2_txdetectrx(iffcq22txdetectrxloopback),
.ch2_txdlyalignerr(iffcq22txdelayalignerr),
.ch2_txdlyalignreq(iffcq22txdelayalignreq),
.ch2_txmldchaindone(iffcq22txmldchaindone),
.ch2_txpcsresetmask(iffcq22txpcsresetmask),
.ch2_txpicodereset(iffcq22txtxpicodereset),
.ch2_txpmaresetdone(iffcq22txpmaresetdone),
.ch2_txpmaresetmask(iffcq22txpmaresetmask),
.ch2_txprbsforceerr(iffcq22txprbsforceerr),
.ch2_txprogdivreset(iffcq22txprogdivreset),
.ch2_txswingouthigh(iffcq22txswingouthigh),
.ch2_rxphaligndone(iffcq22rxphasealigndone),
.ch2_txphaligndone(iffcq22txphasealigndone),
.ch2_rxbyteisaligned(iffcq22rxbyteisaligned),
.ch2_rxdapicodereset(iffcq22rxdapicodereset),
.ch2_rxdapiresetdone(iffcq22rxdapiresetdone),
.ch2_rxdapiresetmask(iffcq22rxdapiresetmask),
.ch2_rxfinealigndone(iffcq22rxfinealigndone),
.ch2_rxphshift180(iffcq22rxphaseshift180req),
.ch2_txdapicodereset(iffcq22txdapicodereset),
.ch2_txdapiresetdone(iffcq22txdapiresetdone),
.ch2_txdapiresetmask(iffcq22txdapiresetmask),
.ch2_txphalignoutrsvd(iffcq22txchicooutrsvd),
.ch2_txphshift180(iffcq22txphaseshift180req),
.ch2_txpicodeovrden(iffcq22txtxpicodeovrden),
.ch2_rxphsetinitreq(iffcq22rxphasesetinitreq),
.ch2_txphsetinitreq(iffcq22txphasesetinitreq),
.ch2_eyescandataerror(iffcq22eyescandataerror),
.ch2_rxdapicodeovrden(iffcq22rxdapicodeovrden),
.ch2_rxmlfinealignreq(iffcq22rxmlfinealignreq),
.ch2_txdapicodeovrden(iffcq22txdapicodeovrden),
.ch2_rxmstresetdone(iffctrlq2mstrxresetdone[2]),
.ch2_rxphsetinitdone(iffcq22rxphasesetinitdone),
.ch2_txmstresetdone(iffctrlq2msttxresetdone[2]),
.ch2_txphsetinitdone(iffcq22txphasesetinitdone),
.ch2_rxdlyalignprog(iffcq22rxdelayalignprogress),
.ch2_rxphalignresetmask(iffcq22rxchicoresetmask),
.ch2_txdlyalignprog(iffcq22txdelayalignprogress),
.ch2_txpausedelayalign(iffcq22txpausedelayalign),
.ch2_txphalignresetmask(iffcq22txchicoresetmask),
.ch2_xpipe5_pipeline_en(iffcq22xpipe5pipelineen),
.ch2_phyesmadaptsave(iffcq22phyesmadaptationsave),
.ch2_rxphshift180done(iffcq22rxphaseshift180done),
.ch2_tx10gstat(iffcq22txethernetstattxlocalfault),
.ch2_txphshift180done(iffcq22txphaseshift180done),
.ch2_rxprogdivresetdone(iffcq22rxprogdivresetdone),
.ch2_rxsimplexphystatus(iffcq22rxsimplexphystatus),
.ch2_txprogdivresetdone(iffcq22txprogdivresetdone),
.ch2_txsimplexphystatus(iffcq22txsimplexphystatus),
.ch2_rxphdlyresetdone(iffcq22rxphasedelayresetdone),
.ch2_txphdlyresetdone(iffcq22txphasedelayresetdone),

.ch3_rxdata(iffcq23rxdata),
.ch3_rxrate(iffcq23rxrate),
.ch3_txdata(iffcq23txdata),
.ch3_txrate(iffcq23txrate),
.ch3_bufgtce(iffcq23bufgtce),
.ch3_gtrsvd(iffcq23pinrsrvd),
.ch3_pcierstb(iffcq23perstb),
.ch3_rxctrl0(iffcq23rxctrl0),
.ch3_rxctrl1(iffcq23rxctrl1),
.ch3_rxctrl2(iffcq23rxctrl2),
.ch3_rxctrl3(iffcq23rxctrl3),
.ch3_rxlpmen(iffcq23rxlpmen),
.ch3_rxpkdet(q2_ch3_rxpkdet),
.ch3_rxqpien(iffcq23rxqpien),
.ch3_rxslide(iffcq23rxslide),
.ch3_rxvalid(iffcq23rxvalid),
.ch3_tstclk0(iffcq23tstclk0),
.ch3_tstclk1(iffcq23tstclk1),
.ch3_txctrl0(iffcq23txctrl0),
.ch3_txctrl1(iffcq23txctrl1),
.ch3_txctrl2(iffcq23txctrl2),
.ch3_txpippmen(iffcq23enppm),
.ch3_txswing(iffcq23txswing),
.ch3_rxpd(iffcq23rxpowerdown),
.ch3_txpd(iffcq23txpowerdown),
.ch3_bufgtdiv(iffcq23bufgtdiv),
.ch3_bufgtrst(iffcq23bufgtrst),
.ch3_iloreset(iffcq23iloreset),
.ch3_loopback(iffcq23loopback),
.ch3_phyready(iffcq23phyready),
.ch3_rxcdrhold(iffcq23cdrhold),
.ch3_rxcdrlock(iffcq23cdrlock),
.ch3_rxheader(iffcq23rxheader),
.ch3_rxlatclk(iffcq23rxlatclk),
.ch3_rxoutclk(q2_ch3_rxoutclk),
.ch3_rxstatus(iffcq23rxstatus),
.ch3_rxusrclk(iffcq23rxusrclk),
.ch3_txcomsas(iffcq23txcomsas),
.ch3_txdeemph(iffcq23txdeemph),
.ch3_txheader(iffcq23txheader),
.ch3_txlatclk(iffcq23txlatclk),
.ch3_txmargin(iffcq23txmargin),
.ch3_txoutclk(q2_ch3_txoutclk),
.ch3_txusrclk(iffcq23txusrclk),
.ch3_dfehold(iffcq23aptexthold),
.ch3_rxuserrdy(iffcq23rxusrrdy),
.ch3_txuserrdy(iffcq23txusrrdy),
.ch3_cdrfreqos(iffcq23cdrfreqos),
.ch3_cdrstepsq(iffcq23cdrstepsq),
.ch3_cdrstepsx(iffcq23cdrstepsx),
.ch3_dfeovrd(iffcq23aptoverwren),
.ch3_dmonitorclk(iffcq23dmonclk),
.ch3_dmonitorout(iffcq23dmonout),
.ch3_gtrxreset(iffcq23gtrxreset),
.ch3_gttxreset(iffcq23gttxreset),
.ch3_pcsrsvdin(iffcq23pcsrsvdin),
.ch3_phystatus(iffcq23phystatus),
.ch3_rxchbondi(iffcq23rxchbondi),
.ch3_rxchbondo(iffcq23rxchbondo),
.ch3_rxprbserr(iffcq23rxprbserr),
.ch3_rxprbssel(iffcq23rxprbssel),
.ch3_rxqpisenn(iffcq23rxqpisenn),
.ch3_rxqpisenp(iffcq23rxqpisenp),
.ch3_txcominit(iffcq23txcominit),
.ch3_txcomwake(iffcq23txcomwake),
.ch3_txdccdone(iffcq23txdccdone),
.ch3_txdiffctrl(iffcq23txdrvamp),
.ch3_txinhibit(iffcq23txinhibit),
.ch3_txpisopd(iffcq23txserpwrdn),
.ch3_txprbssel(iffcq23txprbssel),
.ch3_txqpisenn(iffcq23txqpisenn),
.ch3_txqpisenp(iffcq23txqpisenp),
.ch3_clkrsvd0(iffcq23ckpinrsrvd0),
.ch3_clkrsvd1(iffcq23ckpinrsrvd1),
.ch3_pinrsvdas(iffcq23pinrsrvdas),
.ch3_rxcdrovrden(iffcq23cdrovren),
.ch3_rxosintdone(iffcq23cfokdone),
.ch3_txprecursor(iffcq23txemppre),
.ch3_cdrstepdir(iffcq23cdrstepdir),
.ch3_pcsrsvdout(iffcq23pcsrsvdout),
.ch3_refdebugout(iffcq23refclkpma),
.ch3_rxcdrreset(iffcq23cdrphreset),
.ch3_rxcommadet(iffcq23rxcommadet),
.ch3_rxcomsasdet(iffcq23comsasdet),
.ch3_rxelecidle(iffcq23rxelecidle),
.ch3_rxoobreset(iffcq23rxoobreset),
.ch3_rxpolarity(iffcq23rxpolarity),
.ch3_rxsliderdy(iffcq23rxsliderdy),
.ch3_rxslipdone(iffcq23rxslipdone),
.ch3_rxsyncdone(iffcq23rxsyncdone),
.ch3_txelecidle(iffcq23txelecidle),
.ch3_txpolarity(iffcq23txpolarity),
.ch3_txpostcursor(iffcq23txemppos),
.ch3_txsequence(iffcq23txsequence),
.ch3_txsyncdone(iffcq23txsyncdone),
.ch3_cdrbmcdrreq(iffcq23cdrbmcdreq),
.ch3_rxclkcorcnt(iffcq23rxckcorcnt),
.ch3_txmaincursor(iffcq23txempmain),
.ch3_bufgtcemask(iffcq23bufgtcemask),
.ch3_cdrincpctrl(iffcq23cdrincpctrl),
.ch3_rxbufstatus(iffcq23rxbufstatus),
.ch3_rxcdrphdone(iffcq23rxcdrphdone),
.ch3_rxcominitdet(iffcq23cominitdet),
.ch3_rxcomwakedet(iffcq23comwakedet),
.ch3_rxdapireset(iffcq23rxdapireset),
.ch3_rxdatavalid(iffcq23rxdatavalid),
.ch3_rxresetdone(iffcq23rxresetdone),
.ch3_rxresetmode(iffcq23rxresetmode),
.ch3_rxsyncallin(iffcq23rxsyncallin),
.ch3_txbufstatus(iffcq23txbufstatus),
.ch3_txcomfinish(iffcq23txcomfinish),
.ch3_txdapireset(iffcq23txdapireset),
.ch3_txoneszeros(iffcq23txoneszeros),
.ch3_txqpibiasen(iffcq23txqpibiasen),
.ch3_txqpiweakpu(iffcq23txqpiweakpu),
.ch3_txresetdone(iffcq23txresetdone),
.ch3_txresetmode(iffcq23txresetmode),
.ch3_txsyncallin(iffcq23txsyncallin),
.ch3_rxphdlypd(iffcq23rxphasealignpd),
.ch3_txphdlypd(iffcq23txphasealignpd),
.ch3_bufgtrstmask(iffcq23bufgtrstmask),
.ch3_eyescanreset(iffcq23eyescanreset),
.ch3_hsdppcsreset(iffcq23hsdppcsreset),
.ch3_iloresetdone(iffcq23iloresetdone),
.ch3_iloresetmask(iffcq23iloresetmask),
.ch3_rxdebugpcsout(iffcq23rxoutpcsclk),
.ch3_rxeqtraining(iffcq23rxeqtraining),
.ch3_rxphdlyreset(iffcq23rxphdlyreset),
.ch3_rxprbslocked(iffcq23rxprbslocked),
.ch3_rxstartofseq(iffcq23rxstartofseq),
.ch3_txdebugpcsout(iffcq23txoutpcsclk),
.ch3_txphdlyreset(iffcq23txphdlyreset),
.ch3_rxmstreset(iffctrlq2mstrxreset[3]),
.ch3_txmstreset(iffctrlq2msttxreset[3]),
.ch3_dmonfiforeset(iffcq23dmonfiforeset),
.ch3_rx10gstat(iffcq23rxethernetstatout),
.ch3_rxbyterealign(q2_ch3_rxbyterealign),
.ch3_rxchanbondseq(iffcq23rxchanbondseq),
.ch3_rxchanrealign(iffcq23rxchanrealign),
.ch3_rxgearboxslip(iffcq23rxgearboxslip),
.ch3_rxheadervalid(iffcq23rxheadervalid),
.ch3_rxmldchainreq(iffcq23rxmldchainreq),
.ch3_rxtermination(iffcq23rxtermination),
.ch3_txmldchainreq(iffcq23txmldchainreq),
.ch3_txpippmstepsize(iffcq23stepsizeppm),
.ch3_txswingoutlow(iffcq23txswingoutlow),
.ch3_rxphalignerr(iffcq23rxphasealignerr),
.ch3_rxphalignreq(iffcq23rxphasealignreq),
.ch3_txphalignerr(iffcq23txphasealignerr),
.ch3_txphalignreq(iffcq23txphasealignreq),
.ch3_txphdlytstclk(iffcq23tcoclkfsmfrout),
.ch3_dmonitoroutclk(q2_ch3_dmonitoroutclk),
.ch3_eyescantrigger(iffcq23eyescantrigger),
.ch3_resetexception(iffcq23resetexception),
.ch3_rxchanisaligned(iffcq23rxchisaligned),
.ch3_rxdlyalignerr(iffcq23rxdelayalignerr),
.ch3_rxdlyalignreq(iffcq23rxdelayalignreq),
.ch3_rxmldchaindone(iffcq23rxmldchaindone),
.ch3_rxpcsresetmask(iffcq23rxpcsresetmask),
.ch3_rxpmaresetdone(iffcq23rxpmaresetdone),
.ch3_rxpmaresetmask(iffcq23rxpmaresetmask),
.ch3_rxprbscntreset(iffcq23rxprbscntreset),
.ch3_rxprogdivreset(iffcq23rxprogdivreset),
.ch3_txdetectrx(iffcq23txdetectrxloopback),
.ch3_txdlyalignerr(iffcq23txdelayalignerr),
.ch3_txdlyalignreq(iffcq23txdelayalignreq),
.ch3_txmldchaindone(iffcq23txmldchaindone),
.ch3_txpcsresetmask(iffcq23txpcsresetmask),
.ch3_txpicodereset(iffcq23txtxpicodereset),
.ch3_txpmaresetdone(iffcq23txpmaresetdone),
.ch3_txpmaresetmask(iffcq23txpmaresetmask),
.ch3_txprbsforceerr(iffcq23txprbsforceerr),
.ch3_txprogdivreset(iffcq23txprogdivreset),
.ch3_txswingouthigh(iffcq23txswingouthigh),
.ch3_rxphaligndone(iffcq23rxphasealigndone),
.ch3_txphaligndone(iffcq23txphasealigndone),
.ch3_rxbyteisaligned(iffcq23rxbyteisaligned),
.ch3_rxdapicodereset(iffcq23rxdapicodereset),
.ch3_rxdapiresetdone(iffcq23rxdapiresetdone),
.ch3_rxdapiresetmask(iffcq23rxdapiresetmask),
.ch3_rxfinealigndone(iffcq23rxfinealigndone),
.ch3_rxphshift180(iffcq23rxphaseshift180req),
.ch3_txdapicodereset(iffcq23txdapicodereset),
.ch3_txdapiresetdone(iffcq23txdapiresetdone),
.ch3_txdapiresetmask(iffcq23txdapiresetmask),
.ch3_txphalignoutrsvd(iffcq23txchicooutrsvd),
.ch3_txphshift180(iffcq23txphaseshift180req),
.ch3_txpicodeovrden(iffcq23txtxpicodeovrden),
.ch3_rxphsetinitreq(iffcq23rxphasesetinitreq),
.ch3_txphsetinitreq(iffcq23txphasesetinitreq),
.ch3_eyescandataerror(iffcq23eyescandataerror),
.ch3_rxdapicodeovrden(iffcq23rxdapicodeovrden),
.ch3_rxmlfinealignreq(iffcq23rxmlfinealignreq),
.ch3_txdapicodeovrden(iffcq23txdapicodeovrden),
.ch3_rxmstresetdone(iffctrlq2mstrxresetdone[3]),
.ch3_rxphsetinitdone(iffcq23rxphasesetinitdone),
.ch3_txmstresetdone(iffctrlq2msttxresetdone[3]),
.ch3_txphsetinitdone(iffcq23txphasesetinitdone),
.ch3_rxdlyalignprog(iffcq23rxdelayalignprogress),
.ch3_rxphalignresetmask(iffcq23rxchicoresetmask),
.ch3_txdlyalignprog(iffcq23txdelayalignprogress),
.ch3_txpausedelayalign(iffcq23txpausedelayalign),
.ch3_txphalignresetmask(iffcq23txchicoresetmask),
.ch3_xpipe5_pipeline_en(iffcq23xpipe5pipelineen),
.ch3_phyesmadaptsave(iffcq23phyesmadaptationsave),
.ch3_rxphshift180done(iffcq23rxphaseshift180done),
.ch3_tx10gstat(iffcq23txethernetstattxlocalfault),
.ch3_txphshift180done(iffcq23txphaseshift180done),
.ch3_rxprogdivresetdone(iffcq23rxprogdivresetdone),
.ch3_rxsimplexphystatus(iffcq23rxsimplexphystatus),
.ch3_txprogdivresetdone(iffcq23txprogdivresetdone),
.ch3_txsimplexphystatus(iffcq23txsimplexphystatus),
.ch3_rxphdlyresetdone(iffcq23rxphasedelayresetdone),
.ch3_txphdlyresetdone(iffcq23txphasedelayresetdone),

.ctrlrsvdin(iffctrlq2gtrsvdin),
.ctrlrsvdout(iffctrlq2gtrsvdout),
.coestatusdebug(iffctrlq2coeregrst),
.correcterr(iffctrlq2correctableerr),

.debugtraceclk(iffctrlq2debugtraceclk),
.debugtracetdata(iffctrlq2debugtracetdata),
.debugtraceready(iffctrlq2debugtracetready),
.debugtracetvalid(iffctrlq2debugtracetvalid),

.gpi(iffctrlq2ubgpi),
.gpo(iffctrlq2ubgpo),
.gtpowergood(iffctrlq2gtpowergood),

.hsclk0_rpllpd(iffhsq20rpllpwrdn),
.hsclk0_lcpllpd(iffhsq20lcpllpwrdn),
.hsclk0_rpllfbdiv(iffhsq20rpllfbdiv),
.hsclk0_rpllreset(iffhsq20rpllreset),
.hsclk0_lcpllfbdiv(iffhsq20lcpllfbdiv),
.hsclk0_lcpllreset(iffhsq20lcpllreset),
.hsclk0_rplllock(iffhsq20rpllfreqlock),
.hsclk0_lcplllock(iffhsq20lcpllfreqlock),
.hsclk0_rpllsdmdata(iffhsq20rpllsdmdata),
.hsclk0_rpllfbclklost(iffhsq20rpllfbloss),
.hsclk0_lcpllsdmdata(iffhsq20lcpllsdmdata),
.hsclk0_rxrecclkout0(iffhsq20rxrecclkout0),
.hsclk0_rxrecclkout1(iffhsq20rxrecclkout1),
.hsclk0_lcpllfbclklost(iffhsq20lcpllfbloss),
.hsclk0_rpllrefclklost(iffhsq20rpllrefloss),
.hsclk0_rpllrefclksel(iffhsq20rpllrefseldyn),
.hsclk0_rpllresetmask(iffhsq20rpllresetmask),
.hsclk0_rpllsdmtoggle(iffhsq20rpllsdmtoggle),
.hsclk0_lcpllrefclklost(iffhsq20lcpllrefloss),
.hsclk0_lcpllrefclksel(iffhsq20lcpllrefseldyn),
.hsclk0_lcpllresetmask(iffhsq20lcpllresetmask),
.hsclk0_lcpllsdmtoggle(iffhsq20lcpllsdmtoggle),
.hsclk0_rpllrefclkmonitor(iffhsq20mgtrpllrefclkfa),
.hsclk0_lcpllrefclkmonitor(iffhsq20mgtlcpllrefclkfa),
.hsclk0_rpllresetbypassmode(iffhsq20rpllresetbypassmode),
.hsclk0_lcpllresetbypassmode(iffhsq20lcpllresetbypassmode),

.hsclk1_rpllpd(iffhsq21rpllpwrdn),
.hsclk1_lcpllpd(iffhsq21lcpllpwrdn),
.hsclk1_rpllfbdiv(iffhsq21rpllfbdiv),
.hsclk1_rpllreset(iffhsq21rpllreset),
.hsclk1_lcpllfbdiv(iffhsq21lcpllfbdiv),
.hsclk1_lcpllreset(iffhsq21lcpllreset),
.hsclk1_rplllock(iffhsq21rpllfreqlock),
.hsclk1_lcplllock(iffhsq21lcpllfreqlock),
.hsclk1_rpllsdmdata(iffhsq21rpllsdmdata),
.hsclk1_rpllfbclklost(iffhsq21rpllfbloss),
.hsclk1_lcpllsdmdata(iffhsq21lcpllsdmdata),
.hsclk1_rxrecclkout0(iffhsq21rxrecclkout0),
.hsclk1_rxrecclkout1(iffhsq21rxrecclkout1),
.hsclk1_lcpllfbclklost(iffhsq21lcpllfbloss),
.hsclk1_rpllrefclklost(iffhsq21rpllrefloss),
.hsclk1_rpllrefclksel(iffhsq21rpllrefseldyn),
.hsclk1_rpllresetmask(iffhsq21rpllresetmask),
.hsclk1_rpllsdmtoggle(iffhsq21rpllsdmtoggle),
.hsclk1_lcpllrefclklost(iffhsq21lcpllrefloss),
.hsclk1_lcpllrefclksel(iffhsq21lcpllrefseldyn),
.hsclk1_lcpllresetmask(iffhsq21lcpllresetmask),
.hsclk1_lcpllsdmtoggle(iffhsq21lcpllsdmtoggle),
.hsclk1_rpllrefclkmonitor(iffhsq21mgtrpllrefclkfa),
.hsclk1_lcpllrefclkmonitor(iffhsq21mgtlcpllrefclkfa),
.hsclk1_rpllresetbypassmode(iffhsq21rpllresetbypassmode),
.hsclk1_lcpllresetbypassmode(iffhsq21lcpllresetbypassmode),

.m0_axis_tdata(iffctrlq2m0axistdata),
.m0_axis_tlast(iffctrlq2m0axistlast),
.m1_axis_tdata(iffctrlq2m1axistdata),
.m1_axis_tlast(iffctrlq2m1axistlast),
.m2_axis_tdata(iffctrlq2m2axistdata),
.m2_axis_tlast(iffctrlq2m2axistlast),
.s0_axis_tdata(iffctrlq2s0axistdata),
.s0_axis_tlast(iffctrlq2s0axistlast),
.s1_axis_tdata(iffctrlq2s1axistdata),
.s1_axis_tlast(iffctrlq2s1axistlast),
.s2_axis_tdata(iffctrlq2s2axistdata),
.s2_axis_tlast(iffctrlq2s2axistlast),
.m0_axis_tready(iffctrlq2m0axistready),
.m0_axis_tvalid(iffctrlq2m0axistvalid),
.m1_axis_tready(iffctrlq2m1axistready),
.m1_axis_tvalid(iffctrlq2m1axistvalid),
.m2_axis_tready(iffctrlq2m2axistready),
.m2_axis_tvalid(iffctrlq2m2axistvalid),
.s0_axis_tready(iffctrlq2s0axistready),
.s0_axis_tvalid(iffctrlq2s0axistvalid),
.s1_axis_tready(iffctrlq2s1axistready),
.s1_axis_tvalid(iffctrlq2s1axistvalid),
.s2_axis_tready(iffctrlq2s2axistready),
.s2_axis_tvalid(iffctrlq2s2axistvalid),

.rcalenb(iffctrlq2rcalenb),
.pcieltssm(iffctrlq2pcieltssmstate),
.uncorrecterr(iffctrlq2uncorrectableerr),
.pcielinkreachtarget(iffctrlq2pcielinkreachtarget),

.refclk0_clktestsigint(),
.refclk1_clktestsigint(),
.refclk0_gtrefclkpd(iffrckq20refclkpd),
.refclk1_gtrefclkpd(iffrckq21refclkpd),
.refclk0_clktestsig(iffrckq20hrowtestck),
.refclk1_clktestsig(iffrckq21hrowtestck),
.refclk0_gtrefclkpdint(gt2_refclk0_pdint),
.refclk1_gtrefclkpdint(gt2_refclk1_pdint),

.rxmarginclk(iffctrlq2rxmarginclk),
.rxmarginreqack(iffctrlq2rxmarginreqack),
.rxmarginreqcmd(iffctrlq2rxmarginreqcmd),
.rxmarginreqreq(iffctrlq2rxmarginreqreq),
.rxmarginresack(iffctrlq2rxmarginresack),
.rxmarginrescmd(iffctrlq2rxmarginrescmd),
.rxmarginresreq(iffctrlq2rxmarginresreq),
.rxmarginrespayld(iffctrlq2rxmarginrespayld),
.rxmarginreqpayld(iffctrlq2rxmarginreqpayload),
.rxmarginreqlanenum(iffctrlq2rxmarginreqlanenum),
.rxmarginreslanenum(iffctrlq2rxmarginreslanenum),

.trigin0(iffctrlq2trigin0),
.trigout0(iffctrlq2trigout0),
.trigackin0(iffctrlq2trigackin0),
.trigackout0(iffctrlq2trigackout0),

.ubintr(iffctrlq2ubintr),
.ubmbrst(iffctrlq2ubmbrst),
.ubenable(iffctrlq2ubenable),
.ubrxuart(iffctrlq2ubrxuart),
.ubtxuart(iffctrlq2ubtxuart),
.ubiolmbrst(iffctrlq2ubiolmbrst),
.ubinterrupt(iffctrlq2ubinterrupt),

.pipenorthin(pipenorthoutq1_to_pipenorthinq2),
.pipenorthout(pipenorthoutq2_to_pipenorthinq3),
.rxpisouthin(rxpisouthin_q2_to_rxpsouthout_q3),
.txpisouthin(txpisouthin_q2_to_txpsouthout_q3),
.pipesouthin(pipesouthin_q2_to_pipesouthout_q3),
.rxpinorthin(rxpinorthout_q1_to_rxpinorthin_q2),
.rxpisouthout(rxpisouthin_q1_to_rxpsouthout_q2),
.txpinorthin(txpinorthout_q1_to_txpinorthin_q2),
.txpisouthout(txpisouthin_q1_to_txpsouthout_q2),
.pipesouthout(pipesouthin_q1_to_pipesouthout_q2),
.rxpinorthout(rxpinorthout_q2_to_rxpinorthin_q3),
.txpinorthout(txpinorthout_q2_to_txpinorthin_q3),
.resetdone_northin(resetdone_northout_q1_to_resetdone_northin_q2),
.resetdone_southin(resetdone_southin_q2_to_resetdone_southout_q3),
.resetdone_northout(resetdone_northout_q2_to_resetdone_northin_q3),
.resetdone_southout(resetdone_southin_q1_to_resetdone_southout_q2),

.rxn(gt2_serial_rxn),
.rxp(gt2_serial_rxp),
.txn(gt2_serial_txn),
.txp(gt2_serial_txp)
