.GT_REFCLK0(gt_refclk0_out),

.apb3clk(iffctrlq1apb3clk),
.axisclk(iffctrlq1axisclk),

.apb3psel(iffctrlq1psel),
.apb3paddr(iffctrlq1paddr),
.apb3prdata(iffctrlq1prdata),
.apb3pready(iffctrlq1pready),
.apb3pwdata(iffctrlq1pwdata),
.apb3pwrite(iffctrlq1pwrite),
.apb3penable(iffctrlq1penable),
.apb3presetn(iffctrlq1presetn),
.apb3pslverr(iffctrlq1pslverr),

.bgpdb(iffctrlq1bgpwrdnb),
.bgbypassb(iffctrlq1bgbypass),
.bgrcalovrd(iffctrlq1bgrcalctl),
.bgmonitorenb(iffctrlq1bgtesten),
.bgrcalovrdenb(iffctrlq1bgrcalovrdenb),

.ch0_rxdata(iffcq10rxdata),
.ch0_rxrate(iffcq10rxrate),
.ch0_txdata(iffcq10txdata),
.ch0_txrate(iffcq10txrate),
.ch0_bufgtce(iffcq10bufgtce),
.ch0_gtrsvd(iffcq10pinrsrvd),
.ch0_pcierstb(iffcq10perstb),
.ch0_rxctrl0(iffcq10rxctrl0),
.ch0_rxctrl1(iffcq10rxctrl1),
.ch0_rxctrl2(iffcq10rxctrl2),
.ch0_rxctrl3(iffcq10rxctrl3),
.ch0_rxlpmen(iffcq10rxlpmen),
.ch0_rxpkdet(q1_ch0_rxpkdet),
.ch0_rxqpien(iffcq10rxqpien),
.ch0_rxslide(iffcq10rxslide),
.ch0_rxvalid(iffcq10rxvalid),
.ch0_tstclk0(iffcq10tstclk0),
.ch0_tstclk1(iffcq10tstclk1),
.ch0_txctrl0(iffcq10txctrl0),
.ch0_txctrl1(iffcq10txctrl1),
.ch0_txctrl2(iffcq10txctrl2),
.ch0_txpippmen(iffcq10enppm),
.ch0_txswing(iffcq10txswing),
.ch0_rxpd(iffcq10rxpowerdown),
.ch0_txpd(iffcq10txpowerdown),
.ch0_bufgtdiv(iffcq10bufgtdiv),
.ch0_bufgtrst(iffcq10bufgtrst),
.ch0_iloreset(iffcq10iloreset),
.ch0_loopback(iffcq10loopback),
.ch0_phyready(iffcq10phyready),
.ch0_rxcdrhold(iffcq10cdrhold),
.ch0_rxcdrlock(iffcq10cdrlock),
.ch0_rxheader(iffcq10rxheader),
.ch0_rxlatclk(iffcq10rxlatclk),
.ch0_rxoutclk(q1_ch0_rxoutclk),
.ch0_rxstatus(iffcq10rxstatus),
.ch0_rxusrclk(iffcq10rxusrclk),
.ch0_txcomsas(iffcq10txcomsas),
.ch0_txdeemph(iffcq10txdeemph),
.ch0_txheader(iffcq10txheader),
.ch0_txlatclk(iffcq10txlatclk),
.ch0_txmargin(iffcq10txmargin),
.ch0_txoutclk(q1_ch0_txoutclk),
.ch0_txusrclk(iffcq10txusrclk),
.ch0_dfehold(iffcq10aptexthold),
.ch0_rxuserrdy(iffcq10rxusrrdy),
.ch0_txuserrdy(iffcq10txusrrdy),
.ch0_cdrfreqos(iffcq10cdrfreqos),
.ch0_cdrstepsq(iffcq10cdrstepsq),
.ch0_cdrstepsx(iffcq10cdrstepsx),
.ch0_dfeovrd(iffcq10aptoverwren),
.ch0_dmonitorclk(iffcq10dmonclk),
.ch0_dmonitorout(iffcq10dmonout),
.ch0_gtrxreset(iffcq10gtrxreset),
.ch0_gttxreset(iffcq10gttxreset),
.ch0_pcsrsvdin(iffcq10pcsrsvdin),
.ch0_phystatus(iffcq10phystatus),
.ch0_rxchbondi(iffcq10rxchbondi),
.ch0_rxchbondo(iffcq10rxchbondo),
.ch0_rxprbserr(iffcq10rxprbserr),
.ch0_rxprbssel(iffcq10rxprbssel),
.ch0_rxqpisenn(iffcq10rxqpisenn),
.ch0_rxqpisenp(iffcq10rxqpisenp),
.ch0_txcominit(iffcq10txcominit),
.ch0_txcomwake(iffcq10txcomwake),
.ch0_txdccdone(iffcq10txdccdone),
.ch0_txdiffctrl(iffcq10txdrvamp),
.ch0_txinhibit(iffcq10txinhibit),
.ch0_txpisopd(iffcq10txserpwrdn),
.ch0_txprbssel(iffcq10txprbssel),
.ch0_txqpisenn(iffcq10txqpisenn),
.ch0_txqpisenp(iffcq10txqpisenp),
.ch0_clkrsvd0(iffcq10ckpinrsrvd0),
.ch0_clkrsvd1(iffcq10ckpinrsrvd1),
.ch0_pinrsvdas(iffcq10pinrsrvdas),
.ch0_rxcdrovrden(iffcq10cdrovren),
.ch0_rxosintdone(iffcq10cfokdone),
.ch0_txprecursor(iffcq10txemppre),
.ch0_cdrstepdir(iffcq10cdrstepdir),
.ch0_pcsrsvdout(iffcq10pcsrsvdout),
.ch0_refdebugout(iffcq10refclkpma),
.ch0_rxcdrreset(iffcq10cdrphreset),
.ch0_rxcommadet(iffcq10rxcommadet),
.ch0_rxcomsasdet(iffcq10comsasdet),
.ch0_rxelecidle(iffcq10rxelecidle),
.ch0_rxoobreset(iffcq10rxoobreset),
.ch0_rxpolarity(iffcq10rxpolarity),
.ch0_rxsliderdy(iffcq10rxsliderdy),
.ch0_rxslipdone(iffcq10rxslipdone),
.ch0_rxsyncdone(iffcq10rxsyncdone),
.ch0_txelecidle(iffcq10txelecidle),
.ch0_txpolarity(iffcq10txpolarity),
.ch0_txpostcursor(iffcq10txemppos),
.ch0_txsequence(iffcq10txsequence),
.ch0_txsyncdone(iffcq10txsyncdone),
.ch0_cdrbmcdrreq(iffcq10cdrbmcdreq),
.ch0_rxclkcorcnt(iffcq10rxckcorcnt),
.ch0_txmaincursor(iffcq10txempmain),
.ch0_bufgtcemask(iffcq10bufgtcemask),
.ch0_cdrincpctrl(iffcq10cdrincpctrl),
.ch0_rxbufstatus(iffcq10rxbufstatus),
.ch0_rxcdrphdone(iffcq10rxcdrphdone),
.ch0_rxcominitdet(iffcq10cominitdet),
.ch0_rxcomwakedet(iffcq10comwakedet),
.ch0_rxdapireset(iffcq10rxdapireset),
.ch0_rxdatavalid(iffcq10rxdatavalid),
.ch0_rxresetdone(iffcq10rxresetdone),
.ch0_rxresetmode(iffcq10rxresetmode),
.ch0_rxsyncallin(iffcq10rxsyncallin),
.ch0_txbufstatus(iffcq10txbufstatus),
.ch0_txcomfinish(iffcq10txcomfinish),
.ch0_txdapireset(iffcq10txdapireset),
.ch0_txoneszeros(iffcq10txoneszeros),
.ch0_txqpibiasen(iffcq10txqpibiasen),
.ch0_txqpiweakpu(iffcq10txqpiweakpu),
.ch0_txresetdone(iffcq10txresetdone),
.ch0_txresetmode(iffcq10txresetmode),
.ch0_txsyncallin(iffcq10txsyncallin),
.ch0_rxphdlypd(iffcq10rxphasealignpd),
.ch0_txphdlypd(iffcq10txphasealignpd),
.ch0_bufgtrstmask(iffcq10bufgtrstmask),
.ch0_eyescanreset(iffcq10eyescanreset),
.ch0_hsdppcsreset(iffcq10hsdppcsreset),
.ch0_iloresetdone(iffcq10iloresetdone),
.ch0_iloresetmask(iffcq10iloresetmask),
.ch0_rxdebugpcsout(iffcq10rxoutpcsclk),
.ch0_rxeqtraining(iffcq10rxeqtraining),
.ch0_rxphdlyreset(iffcq10rxphdlyreset),
.ch0_rxprbslocked(iffcq10rxprbslocked),
.ch0_rxstartofseq(iffcq10rxstartofseq),
.ch0_txdebugpcsout(iffcq10txoutpcsclk),
.ch0_txphdlyreset(iffcq10txphdlyreset),
.ch0_rxmstreset(iffctrlq1mstrxreset[0]),
.ch0_txmstreset(iffctrlq1msttxreset[0]),
.ch0_dmonfiforeset(iffcq10dmonfiforeset),
.ch0_rx10gstat(iffcq10rxethernetstatout),
.ch0_rxbyterealign(q1_ch0_rxbyterealign),
.ch0_rxchanbondseq(iffcq10rxchanbondseq),
.ch0_rxchanrealign(iffcq10rxchanrealign),
.ch0_rxgearboxslip(iffcq10rxgearboxslip),
.ch0_rxheadervalid(iffcq10rxheadervalid),
.ch0_rxmldchainreq(iffcq10rxmldchainreq),
.ch0_rxtermination(iffcq10rxtermination),
.ch0_txmldchainreq(iffcq10txmldchainreq),
.ch0_txpippmstepsize(iffcq10stepsizeppm),
.ch0_txswingoutlow(iffcq10txswingoutlow),
.ch0_rxphalignerr(iffcq10rxphasealignerr),
.ch0_rxphalignreq(iffcq10rxphasealignreq),
.ch0_txphalignerr(iffcq10txphasealignerr),
.ch0_txphalignreq(iffcq10txphasealignreq),
.ch0_txphdlytstclk(iffcq10tcoclkfsmfrout),
.ch0_dmonitoroutclk(q1_ch0_dmonitoroutclk),
.ch0_eyescantrigger(iffcq10eyescantrigger),
.ch0_resetexception(iffcq10resetexception),
.ch0_rxchanisaligned(iffcq10rxchisaligned),
.ch0_rxdlyalignerr(iffcq10rxdelayalignerr),
.ch0_rxdlyalignreq(iffcq10rxdelayalignreq),
.ch0_rxmldchaindone(iffcq10rxmldchaindone),
.ch0_rxpcsresetmask(iffcq10rxpcsresetmask),
.ch0_rxpmaresetdone(iffcq10rxpmaresetdone),
.ch0_rxpmaresetmask(iffcq10rxpmaresetmask),
.ch0_rxprbscntreset(iffcq10rxprbscntreset),
.ch0_rxprogdivreset(iffcq10rxprogdivreset),
.ch0_txdetectrx(iffcq10txdetectrxloopback),
.ch0_txdlyalignerr(iffcq10txdelayalignerr),
.ch0_txdlyalignreq(iffcq10txdelayalignreq),
.ch0_txmldchaindone(iffcq10txmldchaindone),
.ch0_txpcsresetmask(iffcq10txpcsresetmask),
.ch0_txpicodereset(iffcq10txtxpicodereset),
.ch0_txpmaresetdone(iffcq10txpmaresetdone),
.ch0_txpmaresetmask(iffcq10txpmaresetmask),
.ch0_txprbsforceerr(iffcq10txprbsforceerr),
.ch0_txprogdivreset(iffcq10txprogdivreset),
.ch0_txswingouthigh(iffcq10txswingouthigh),
.ch0_rxphaligndone(iffcq10rxphasealigndone),
.ch0_txphaligndone(iffcq10txphasealigndone),
.ch0_rxbyteisaligned(iffcq10rxbyteisaligned),
.ch0_rxdapicodereset(iffcq10rxdapicodereset),
.ch0_rxdapiresetdone(iffcq10rxdapiresetdone),
.ch0_rxdapiresetmask(iffcq10rxdapiresetmask),
.ch0_rxfinealigndone(iffcq10rxfinealigndone),
.ch0_rxphshift180(iffcq10rxphaseshift180req),
.ch0_txdapicodereset(iffcq10txdapicodereset),
.ch0_txdapiresetdone(iffcq10txdapiresetdone),
.ch0_txdapiresetmask(iffcq10txdapiresetmask),
.ch0_txphalignoutrsvd(iffcq10txchicooutrsvd),
.ch0_txphshift180(iffcq10txphaseshift180req),
.ch0_txpicodeovrden(iffcq10txtxpicodeovrden),
.ch0_rxphsetinitreq(iffcq10rxphasesetinitreq),
.ch0_txphsetinitreq(iffcq10txphasesetinitreq),
.ch0_eyescandataerror(iffcq10eyescandataerror),
.ch0_rxdapicodeovrden(iffcq10rxdapicodeovrden),
.ch0_rxmlfinealignreq(iffcq10rxmlfinealignreq),
.ch0_txdapicodeovrden(iffcq10txdapicodeovrden),
.ch0_rxmstresetdone(iffctrlq1mstrxresetdone[0]),
.ch0_rxphsetinitdone(iffcq10rxphasesetinitdone),
.ch0_txmstresetdone(iffctrlq1msttxresetdone[0]),
.ch0_txphsetinitdone(iffcq10txphasesetinitdone),
.ch0_rxdlyalignprog(iffcq10rxdelayalignprogress),
.ch0_rxphalignresetmask(iffcq10rxchicoresetmask),
.ch0_txdlyalignprog(iffcq10txdelayalignprogress),
.ch0_txpausedelayalign(iffcq10txpausedelayalign),
.ch0_txphalignresetmask(iffcq10txchicoresetmask),
.ch0_xpipe5_pipeline_en(iffcq10xpipe5pipelineen),
.ch0_phyesmadaptsave(iffcq10phyesmadaptationsave),
.ch0_rxphshift180done(iffcq10rxphaseshift180done),
.ch0_tx10gstat(iffcq10txethernetstattxlocalfault),
.ch0_txphshift180done(iffcq10txphaseshift180done),
.ch0_rxprogdivresetdone(iffcq10rxprogdivresetdone),
.ch0_rxsimplexphystatus(iffcq10rxsimplexphystatus),
.ch0_txprogdivresetdone(iffcq10txprogdivresetdone),
.ch0_txsimplexphystatus(iffcq10txsimplexphystatus),
.ch0_rxphdlyresetdone(iffcq10rxphasedelayresetdone),
.ch0_txphdlyresetdone(iffcq10txphasedelayresetdone),

.ch1_rxdata(iffcq11rxdata),
.ch1_rxrate(iffcq11rxrate),
.ch1_txdata(iffcq11txdata),
.ch1_txrate(iffcq11txrate),
.ch1_bufgtce(iffcq11bufgtce),
.ch1_gtrsvd(iffcq11pinrsrvd),
.ch1_pcierstb(iffcq11perstb),
.ch1_rxctrl0(iffcq11rxctrl0),
.ch1_rxctrl1(iffcq11rxctrl1),
.ch1_rxctrl2(iffcq11rxctrl2),
.ch1_rxctrl3(iffcq11rxctrl3),
.ch1_rxlpmen(iffcq11rxlpmen),
.ch1_rxpkdet(q1_ch1_rxpkdet),
.ch1_rxqpien(iffcq11rxqpien),
.ch1_rxslide(iffcq11rxslide),
.ch1_rxvalid(iffcq11rxvalid),
.ch1_tstclk0(iffcq11tstclk0),
.ch1_tstclk1(iffcq11tstclk1),
.ch1_txctrl0(iffcq11txctrl0),
.ch1_txctrl1(iffcq11txctrl1),
.ch1_txctrl2(iffcq11txctrl2),
.ch1_txpippmen(iffcq11enppm),
.ch1_txswing(iffcq11txswing),
.ch1_rxpd(iffcq11rxpowerdown),
.ch1_txpd(iffcq11txpowerdown),
.ch1_bufgtdiv(iffcq11bufgtdiv),
.ch1_bufgtrst(iffcq11bufgtrst),
.ch1_iloreset(iffcq11iloreset),
.ch1_loopback(iffcq11loopback),
.ch1_phyready(iffcq11phyready),
.ch1_rxcdrhold(iffcq11cdrhold),
.ch1_rxcdrlock(iffcq11cdrlock),
.ch1_rxheader(iffcq11rxheader),
.ch1_rxlatclk(iffcq11rxlatclk),
.ch1_rxoutclk(q1_ch1_rxoutclk),
.ch1_rxstatus(iffcq11rxstatus),
.ch1_rxusrclk(iffcq11rxusrclk),
.ch1_txcomsas(iffcq11txcomsas),
.ch1_txdeemph(iffcq11txdeemph),
.ch1_txheader(iffcq11txheader),
.ch1_txlatclk(iffcq11txlatclk),
.ch1_txmargin(iffcq11txmargin),
.ch1_txoutclk(q1_ch1_txoutclk),
.ch1_txusrclk(iffcq11txusrclk),
.ch1_dfehold(iffcq11aptexthold),
.ch1_rxuserrdy(iffcq11rxusrrdy),
.ch1_txuserrdy(iffcq11txusrrdy),
.ch1_cdrfreqos(iffcq11cdrfreqos),
.ch1_cdrstepsq(iffcq11cdrstepsq),
.ch1_cdrstepsx(iffcq11cdrstepsx),
.ch1_dfeovrd(iffcq11aptoverwren),
.ch1_dmonitorclk(iffcq11dmonclk),
.ch1_dmonitorout(iffcq11dmonout),
.ch1_gtrxreset(iffcq11gtrxreset),
.ch1_gttxreset(iffcq11gttxreset),
.ch1_pcsrsvdin(iffcq11pcsrsvdin),
.ch1_phystatus(iffcq11phystatus),
.ch1_rxchbondi(iffcq11rxchbondi),
.ch1_rxchbondo(iffcq11rxchbondo),
.ch1_rxprbserr(iffcq11rxprbserr),
.ch1_rxprbssel(iffcq11rxprbssel),
.ch1_rxqpisenn(iffcq11rxqpisenn),
.ch1_rxqpisenp(iffcq11rxqpisenp),
.ch1_txcominit(iffcq11txcominit),
.ch1_txcomwake(iffcq11txcomwake),
.ch1_txdccdone(iffcq11txdccdone),
.ch1_txdiffctrl(iffcq11txdrvamp),
.ch1_txinhibit(iffcq11txinhibit),
.ch1_txpisopd(iffcq11txserpwrdn),
.ch1_txprbssel(iffcq11txprbssel),
.ch1_txqpisenn(iffcq11txqpisenn),
.ch1_txqpisenp(iffcq11txqpisenp),
.ch1_clkrsvd0(iffcq11ckpinrsrvd0),
.ch1_clkrsvd1(iffcq11ckpinrsrvd1),
.ch1_pinrsvdas(iffcq11pinrsrvdas),
.ch1_rxcdrovrden(iffcq11cdrovren),
.ch1_rxosintdone(iffcq11cfokdone),
.ch1_txprecursor(iffcq11txemppre),
.ch1_cdrstepdir(iffcq11cdrstepdir),
.ch1_pcsrsvdout(iffcq11pcsrsvdout),
.ch1_refdebugout(iffcq11refclkpma),
.ch1_rxcdrreset(iffcq11cdrphreset),
.ch1_rxcommadet(iffcq11rxcommadet),
.ch1_rxcomsasdet(iffcq11comsasdet),
.ch1_rxelecidle(iffcq11rxelecidle),
.ch1_rxoobreset(iffcq11rxoobreset),
.ch1_rxpolarity(iffcq11rxpolarity),
.ch1_rxsliderdy(iffcq11rxsliderdy),
.ch1_rxslipdone(iffcq11rxslipdone),
.ch1_rxsyncdone(iffcq11rxsyncdone),
.ch1_txelecidle(iffcq11txelecidle),
.ch1_txpolarity(iffcq11txpolarity),
.ch1_txpostcursor(iffcq11txemppos),
.ch1_txsequence(iffcq11txsequence),
.ch1_txsyncdone(iffcq11txsyncdone),
.ch1_cdrbmcdrreq(iffcq11cdrbmcdreq),
.ch1_rxclkcorcnt(iffcq11rxckcorcnt),
.ch1_txmaincursor(iffcq11txempmain),
.ch1_bufgtcemask(iffcq11bufgtcemask),
.ch1_cdrincpctrl(iffcq11cdrincpctrl),
.ch1_rxbufstatus(iffcq11rxbufstatus),
.ch1_rxcdrphdone(iffcq11rxcdrphdone),
.ch1_rxcominitdet(iffcq11cominitdet),
.ch1_rxcomwakedet(iffcq11comwakedet),
.ch1_rxdapireset(iffcq11rxdapireset),
.ch1_rxdatavalid(iffcq11rxdatavalid),
.ch1_rxresetdone(iffcq11rxresetdone),
.ch1_rxresetmode(iffcq11rxresetmode),
.ch1_rxsyncallin(iffcq11rxsyncallin),
.ch1_txbufstatus(iffcq11txbufstatus),
.ch1_txcomfinish(iffcq11txcomfinish),
.ch1_txdapireset(iffcq11txdapireset),
.ch1_txoneszeros(iffcq11txoneszeros),
.ch1_txqpibiasen(iffcq11txqpibiasen),
.ch1_txqpiweakpu(iffcq11txqpiweakpu),
.ch1_txresetdone(iffcq11txresetdone),
.ch1_txresetmode(iffcq11txresetmode),
.ch1_txsyncallin(iffcq11txsyncallin),
.ch1_rxphdlypd(iffcq11rxphasealignpd),
.ch1_txphdlypd(iffcq11txphasealignpd),
.ch1_bufgtrstmask(iffcq11bufgtrstmask),
.ch1_eyescanreset(iffcq11eyescanreset),
.ch1_hsdppcsreset(iffcq11hsdppcsreset),
.ch1_iloresetdone(iffcq11iloresetdone),
.ch1_iloresetmask(iffcq11iloresetmask),
.ch1_rxdebugpcsout(iffcq11rxoutpcsclk),
.ch1_rxeqtraining(iffcq11rxeqtraining),
.ch1_rxphdlyreset(iffcq11rxphdlyreset),
.ch1_rxprbslocked(iffcq11rxprbslocked),
.ch1_rxstartofseq(iffcq11rxstartofseq),
.ch1_txdebugpcsout(iffcq11txoutpcsclk),
.ch1_txphdlyreset(iffcq11txphdlyreset),
.ch1_rxmstreset(iffctrlq1mstrxreset[1]),
.ch1_txmstreset(iffctrlq1msttxreset[1]),
.ch1_dmonfiforeset(iffcq11dmonfiforeset),
.ch1_rx10gstat(iffcq11rxethernetstatout),
.ch1_rxbyterealign(q1_ch1_rxbyterealign),
.ch1_rxchanbondseq(iffcq11rxchanbondseq),
.ch1_rxchanrealign(iffcq11rxchanrealign),
.ch1_rxgearboxslip(iffcq11rxgearboxslip),
.ch1_rxheadervalid(iffcq11rxheadervalid),
.ch1_rxmldchainreq(iffcq11rxmldchainreq),
.ch1_rxtermination(iffcq11rxtermination),
.ch1_txmldchainreq(iffcq11txmldchainreq),
.ch1_txpippmstepsize(iffcq11stepsizeppm),
.ch1_txswingoutlow(iffcq11txswingoutlow),
.ch1_rxphalignerr(iffcq11rxphasealignerr),
.ch1_rxphalignreq(iffcq11rxphasealignreq),
.ch1_txphalignerr(iffcq11txphasealignerr),
.ch1_txphalignreq(iffcq11txphasealignreq),
.ch1_txphdlytstclk(iffcq11tcoclkfsmfrout),
.ch1_dmonitoroutclk(q1_ch1_dmonitoroutclk),
.ch1_eyescantrigger(iffcq11eyescantrigger),
.ch1_resetexception(iffcq11resetexception),
.ch1_rxchanisaligned(iffcq11rxchisaligned),
.ch1_rxdlyalignerr(iffcq11rxdelayalignerr),
.ch1_rxdlyalignreq(iffcq11rxdelayalignreq),
.ch1_rxmldchaindone(iffcq11rxmldchaindone),
.ch1_rxpcsresetmask(iffcq11rxpcsresetmask),
.ch1_rxpmaresetdone(iffcq11rxpmaresetdone),
.ch1_rxpmaresetmask(iffcq11rxpmaresetmask),
.ch1_rxprbscntreset(iffcq11rxprbscntreset),
.ch1_rxprogdivreset(iffcq11rxprogdivreset),
.ch1_txdetectrx(iffcq11txdetectrxloopback),
.ch1_txdlyalignerr(iffcq11txdelayalignerr),
.ch1_txdlyalignreq(iffcq11txdelayalignreq),
.ch1_txmldchaindone(iffcq11txmldchaindone),
.ch1_txpcsresetmask(iffcq11txpcsresetmask),
.ch1_txpicodereset(iffcq11txtxpicodereset),
.ch1_txpmaresetdone(iffcq11txpmaresetdone),
.ch1_txpmaresetmask(iffcq11txpmaresetmask),
.ch1_txprbsforceerr(iffcq11txprbsforceerr),
.ch1_txprogdivreset(iffcq11txprogdivreset),
.ch1_txswingouthigh(iffcq11txswingouthigh),
.ch1_rxphaligndone(iffcq11rxphasealigndone),
.ch1_txphaligndone(iffcq11txphasealigndone),
.ch1_rxbyteisaligned(iffcq11rxbyteisaligned),
.ch1_rxdapicodereset(iffcq11rxdapicodereset),
.ch1_rxdapiresetdone(iffcq11rxdapiresetdone),
.ch1_rxdapiresetmask(iffcq11rxdapiresetmask),
.ch1_rxfinealigndone(iffcq11rxfinealigndone),
.ch1_rxphshift180(iffcq11rxphaseshift180req),
.ch1_txdapicodereset(iffcq11txdapicodereset),
.ch1_txdapiresetdone(iffcq11txdapiresetdone),
.ch1_txdapiresetmask(iffcq11txdapiresetmask),
.ch1_txphalignoutrsvd(iffcq11txchicooutrsvd),
.ch1_txphshift180(iffcq11txphaseshift180req),
.ch1_txpicodeovrden(iffcq11txtxpicodeovrden),
.ch1_rxphsetinitreq(iffcq11rxphasesetinitreq),
.ch1_txphsetinitreq(iffcq11txphasesetinitreq),
.ch1_eyescandataerror(iffcq11eyescandataerror),
.ch1_rxdapicodeovrden(iffcq11rxdapicodeovrden),
.ch1_rxmlfinealignreq(iffcq11rxmlfinealignreq),
.ch1_txdapicodeovrden(iffcq11txdapicodeovrden),
.ch1_rxmstresetdone(iffctrlq1mstrxresetdone[1]),
.ch1_rxphsetinitdone(iffcq11rxphasesetinitdone),
.ch1_txmstresetdone(iffctrlq1msttxresetdone[1]),
.ch1_txphsetinitdone(iffcq11txphasesetinitdone),
.ch1_rxdlyalignprog(iffcq11rxdelayalignprogress),
.ch1_rxphalignresetmask(iffcq11rxchicoresetmask),
.ch1_txdlyalignprog(iffcq11txdelayalignprogress),
.ch1_txpausedelayalign(iffcq11txpausedelayalign),
.ch1_txphalignresetmask(iffcq11txchicoresetmask),
.ch1_xpipe5_pipeline_en(iffcq11xpipe5pipelineen),
.ch1_phyesmadaptsave(iffcq11phyesmadaptationsave),
.ch1_rxphshift180done(iffcq11rxphaseshift180done),
.ch1_tx10gstat(iffcq11txethernetstattxlocalfault),
.ch1_txphshift180done(iffcq11txphaseshift180done),
.ch1_rxprogdivresetdone(iffcq11rxprogdivresetdone),
.ch1_rxsimplexphystatus(iffcq11rxsimplexphystatus),
.ch1_txprogdivresetdone(iffcq11txprogdivresetdone),
.ch1_txsimplexphystatus(iffcq11txsimplexphystatus),
.ch1_rxphdlyresetdone(iffcq11rxphasedelayresetdone),
.ch1_txphdlyresetdone(iffcq11txphasedelayresetdone),

.ch2_rxdata(iffcq12rxdata),
.ch2_rxrate(iffcq12rxrate),
.ch2_txdata(iffcq12txdata),
.ch2_txrate(iffcq12txrate),
.ch2_bufgtce(iffcq12bufgtce),
.ch2_gtrsvd(iffcq12pinrsrvd),
.ch2_pcierstb(iffcq12perstb),
.ch2_rxctrl0(iffcq12rxctrl0),
.ch2_rxctrl1(iffcq12rxctrl1),
.ch2_rxctrl2(iffcq12rxctrl2),
.ch2_rxctrl3(iffcq12rxctrl3),
.ch2_rxlpmen(iffcq12rxlpmen),
.ch2_rxpkdet(q1_ch2_rxpkdet),
.ch2_rxqpien(iffcq12rxqpien),
.ch2_rxslide(iffcq12rxslide),
.ch2_rxvalid(iffcq12rxvalid),
.ch2_tstclk0(iffcq12tstclk0),
.ch2_tstclk1(iffcq12tstclk1),
.ch2_txctrl0(iffcq12txctrl0),
.ch2_txctrl1(iffcq12txctrl1),
.ch2_txctrl2(iffcq12txctrl2),
.ch2_txpippmen(iffcq12enppm),
.ch2_txswing(iffcq12txswing),
.ch2_rxpd(iffcq12rxpowerdown),
.ch2_txpd(iffcq12txpowerdown),
.ch2_bufgtdiv(iffcq12bufgtdiv),
.ch2_bufgtrst(iffcq12bufgtrst),
.ch2_iloreset(iffcq12iloreset),
.ch2_loopback(iffcq12loopback),
.ch2_phyready(iffcq12phyready),
.ch2_rxcdrhold(iffcq12cdrhold),
.ch2_rxcdrlock(iffcq12cdrlock),
.ch2_rxheader(iffcq12rxheader),
.ch2_rxlatclk(iffcq12rxlatclk),
.ch2_rxoutclk(q1_ch2_rxoutclk),
.ch2_rxstatus(iffcq12rxstatus),
.ch2_rxusrclk(iffcq12rxusrclk),
.ch2_txcomsas(iffcq12txcomsas),
.ch2_txdeemph(iffcq12txdeemph),
.ch2_txheader(iffcq12txheader),
.ch2_txlatclk(iffcq12txlatclk),
.ch2_txmargin(iffcq12txmargin),
.ch2_txoutclk(q1_ch2_txoutclk),
.ch2_txusrclk(iffcq12txusrclk),
.ch2_dfehold(iffcq12aptexthold),
.ch2_rxuserrdy(iffcq12rxusrrdy),
.ch2_txuserrdy(iffcq12txusrrdy),
.ch2_cdrfreqos(iffcq12cdrfreqos),
.ch2_cdrstepsq(iffcq12cdrstepsq),
.ch2_cdrstepsx(iffcq12cdrstepsx),
.ch2_dfeovrd(iffcq12aptoverwren),
.ch2_dmonitorclk(iffcq12dmonclk),
.ch2_dmonitorout(iffcq12dmonout),
.ch2_gtrxreset(iffcq12gtrxreset),
.ch2_gttxreset(iffcq12gttxreset),
.ch2_pcsrsvdin(iffcq12pcsrsvdin),
.ch2_phystatus(iffcq12phystatus),
.ch2_rxchbondi(iffcq12rxchbondi),
.ch2_rxchbondo(iffcq12rxchbondo),
.ch2_rxprbserr(iffcq12rxprbserr),
.ch2_rxprbssel(iffcq12rxprbssel),
.ch2_rxqpisenn(iffcq12rxqpisenn),
.ch2_rxqpisenp(iffcq12rxqpisenp),
.ch2_txcominit(iffcq12txcominit),
.ch2_txcomwake(iffcq12txcomwake),
.ch2_txdccdone(iffcq12txdccdone),
.ch2_txdiffctrl(iffcq12txdrvamp),
.ch2_txinhibit(iffcq12txinhibit),
.ch2_txpisopd(iffcq12txserpwrdn),
.ch2_txprbssel(iffcq12txprbssel),
.ch2_txqpisenn(iffcq12txqpisenn),
.ch2_txqpisenp(iffcq12txqpisenp),
.ch2_clkrsvd0(iffcq12ckpinrsrvd0),
.ch2_clkrsvd1(iffcq12ckpinrsrvd1),
.ch2_pinrsvdas(iffcq12pinrsrvdas),
.ch2_rxcdrovrden(iffcq12cdrovren),
.ch2_rxosintdone(iffcq12cfokdone),
.ch2_txprecursor(iffcq12txemppre),
.ch2_cdrstepdir(iffcq12cdrstepdir),
.ch2_pcsrsvdout(iffcq12pcsrsvdout),
.ch2_refdebugout(iffcq12refclkpma),
.ch2_rxcdrreset(iffcq12cdrphreset),
.ch2_rxcommadet(iffcq12rxcommadet),
.ch2_rxcomsasdet(iffcq12comsasdet),
.ch2_rxelecidle(iffcq12rxelecidle),
.ch2_rxoobreset(iffcq12rxoobreset),
.ch2_rxpolarity(iffcq12rxpolarity),
.ch2_rxsliderdy(iffcq12rxsliderdy),
.ch2_rxslipdone(iffcq12rxslipdone),
.ch2_rxsyncdone(iffcq12rxsyncdone),
.ch2_txelecidle(iffcq12txelecidle),
.ch2_txpolarity(iffcq12txpolarity),
.ch2_txpostcursor(iffcq12txemppos),
.ch2_txsequence(iffcq12txsequence),
.ch2_txsyncdone(iffcq12txsyncdone),
.ch2_cdrbmcdrreq(iffcq12cdrbmcdreq),
.ch2_rxclkcorcnt(iffcq12rxckcorcnt),
.ch2_txmaincursor(iffcq12txempmain),
.ch2_bufgtcemask(iffcq12bufgtcemask),
.ch2_cdrincpctrl(iffcq12cdrincpctrl),
.ch2_rxbufstatus(iffcq12rxbufstatus),
.ch2_rxcdrphdone(iffcq12rxcdrphdone),
.ch2_rxcominitdet(iffcq12cominitdet),
.ch2_rxcomwakedet(iffcq12comwakedet),
.ch2_rxdapireset(iffcq12rxdapireset),
.ch2_rxdatavalid(iffcq12rxdatavalid),
.ch2_rxresetdone(iffcq12rxresetdone),
.ch2_rxresetmode(iffcq12rxresetmode),
.ch2_rxsyncallin(iffcq12rxsyncallin),
.ch2_txbufstatus(iffcq12txbufstatus),
.ch2_txcomfinish(iffcq12txcomfinish),
.ch2_txdapireset(iffcq12txdapireset),
.ch2_txoneszeros(iffcq12txoneszeros),
.ch2_txqpibiasen(iffcq12txqpibiasen),
.ch2_txqpiweakpu(iffcq12txqpiweakpu),
.ch2_txresetdone(iffcq12txresetdone),
.ch2_txresetmode(iffcq12txresetmode),
.ch2_txsyncallin(iffcq12txsyncallin),
.ch2_rxphdlypd(iffcq12rxphasealignpd),
.ch2_txphdlypd(iffcq12txphasealignpd),
.ch2_bufgtrstmask(iffcq12bufgtrstmask),
.ch2_eyescanreset(iffcq12eyescanreset),
.ch2_hsdppcsreset(iffcq12hsdppcsreset),
.ch2_iloresetdone(iffcq12iloresetdone),
.ch2_iloresetmask(iffcq12iloresetmask),
.ch2_rxdebugpcsout(iffcq12rxoutpcsclk),
.ch2_rxeqtraining(iffcq12rxeqtraining),
.ch2_rxphdlyreset(iffcq12rxphdlyreset),
.ch2_rxprbslocked(iffcq12rxprbslocked),
.ch2_rxstartofseq(iffcq12rxstartofseq),
.ch2_txdebugpcsout(iffcq12txoutpcsclk),
.ch2_txphdlyreset(iffcq12txphdlyreset),
.ch2_rxmstreset(iffctrlq1mstrxreset[2]),
.ch2_txmstreset(iffctrlq1msttxreset[2]),
.ch2_dmonfiforeset(iffcq12dmonfiforeset),
.ch2_rx10gstat(iffcq12rxethernetstatout),
.ch2_rxbyterealign(q1_ch2_rxbyterealign),
.ch2_rxchanbondseq(iffcq12rxchanbondseq),
.ch2_rxchanrealign(iffcq12rxchanrealign),
.ch2_rxgearboxslip(iffcq12rxgearboxslip),
.ch2_rxheadervalid(iffcq12rxheadervalid),
.ch2_rxmldchainreq(iffcq12rxmldchainreq),
.ch2_rxtermination(iffcq12rxtermination),
.ch2_txmldchainreq(iffcq12txmldchainreq),
.ch2_txpippmstepsize(iffcq12stepsizeppm),
.ch2_txswingoutlow(iffcq12txswingoutlow),
.ch2_rxphalignerr(iffcq12rxphasealignerr),
.ch2_rxphalignreq(iffcq12rxphasealignreq),
.ch2_txphalignerr(iffcq12txphasealignerr),
.ch2_txphalignreq(iffcq12txphasealignreq),
.ch2_txphdlytstclk(iffcq12tcoclkfsmfrout),
.ch2_dmonitoroutclk(q1_ch2_dmonitoroutclk),
.ch2_eyescantrigger(iffcq12eyescantrigger),
.ch2_resetexception(iffcq12resetexception),
.ch2_rxchanisaligned(iffcq12rxchisaligned),
.ch2_rxdlyalignerr(iffcq12rxdelayalignerr),
.ch2_rxdlyalignreq(iffcq12rxdelayalignreq),
.ch2_rxmldchaindone(iffcq12rxmldchaindone),
.ch2_rxpcsresetmask(iffcq12rxpcsresetmask),
.ch2_rxpmaresetdone(iffcq12rxpmaresetdone),
.ch2_rxpmaresetmask(iffcq12rxpmaresetmask),
.ch2_rxprbscntreset(iffcq12rxprbscntreset),
.ch2_rxprogdivreset(iffcq12rxprogdivreset),
.ch2_txdetectrx(iffcq12txdetectrxloopback),
.ch2_txdlyalignerr(iffcq12txdelayalignerr),
.ch2_txdlyalignreq(iffcq12txdelayalignreq),
.ch2_txmldchaindone(iffcq12txmldchaindone),
.ch2_txpcsresetmask(iffcq12txpcsresetmask),
.ch2_txpicodereset(iffcq12txtxpicodereset),
.ch2_txpmaresetdone(iffcq12txpmaresetdone),
.ch2_txpmaresetmask(iffcq12txpmaresetmask),
.ch2_txprbsforceerr(iffcq12txprbsforceerr),
.ch2_txprogdivreset(iffcq12txprogdivreset),
.ch2_txswingouthigh(iffcq12txswingouthigh),
.ch2_rxphaligndone(iffcq12rxphasealigndone),
.ch2_txphaligndone(iffcq12txphasealigndone),
.ch2_rxbyteisaligned(iffcq12rxbyteisaligned),
.ch2_rxdapicodereset(iffcq12rxdapicodereset),
.ch2_rxdapiresetdone(iffcq12rxdapiresetdone),
.ch2_rxdapiresetmask(iffcq12rxdapiresetmask),
.ch2_rxfinealigndone(iffcq12rxfinealigndone),
.ch2_rxphshift180(iffcq12rxphaseshift180req),
.ch2_txdapicodereset(iffcq12txdapicodereset),
.ch2_txdapiresetdone(iffcq12txdapiresetdone),
.ch2_txdapiresetmask(iffcq12txdapiresetmask),
.ch2_txphalignoutrsvd(iffcq12txchicooutrsvd),
.ch2_txphshift180(iffcq12txphaseshift180req),
.ch2_txpicodeovrden(iffcq12txtxpicodeovrden),
.ch2_rxphsetinitreq(iffcq12rxphasesetinitreq),
.ch2_txphsetinitreq(iffcq12txphasesetinitreq),
.ch2_eyescandataerror(iffcq12eyescandataerror),
.ch2_rxdapicodeovrden(iffcq12rxdapicodeovrden),
.ch2_rxmlfinealignreq(iffcq12rxmlfinealignreq),
.ch2_txdapicodeovrden(iffcq12txdapicodeovrden),
.ch2_rxmstresetdone(iffctrlq1mstrxresetdone[2]),
.ch2_rxphsetinitdone(iffcq12rxphasesetinitdone),
.ch2_txmstresetdone(iffctrlq1msttxresetdone[2]),
.ch2_txphsetinitdone(iffcq12txphasesetinitdone),
.ch2_rxdlyalignprog(iffcq12rxdelayalignprogress),
.ch2_rxphalignresetmask(iffcq12rxchicoresetmask),
.ch2_txdlyalignprog(iffcq12txdelayalignprogress),
.ch2_txpausedelayalign(iffcq12txpausedelayalign),
.ch2_txphalignresetmask(iffcq12txchicoresetmask),
.ch2_xpipe5_pipeline_en(iffcq12xpipe5pipelineen),
.ch2_phyesmadaptsave(iffcq12phyesmadaptationsave),
.ch2_rxphshift180done(iffcq12rxphaseshift180done),
.ch2_tx10gstat(iffcq12txethernetstattxlocalfault),
.ch2_txphshift180done(iffcq12txphaseshift180done),
.ch2_rxprogdivresetdone(iffcq12rxprogdivresetdone),
.ch2_rxsimplexphystatus(iffcq12rxsimplexphystatus),
.ch2_txprogdivresetdone(iffcq12txprogdivresetdone),
.ch2_txsimplexphystatus(iffcq12txsimplexphystatus),
.ch2_rxphdlyresetdone(iffcq12rxphasedelayresetdone),
.ch2_txphdlyresetdone(iffcq12txphasedelayresetdone),

.ch3_rxdata(iffcq13rxdata),
.ch3_rxrate(iffcq13rxrate),
.ch3_txdata(iffcq13txdata),
.ch3_txrate(iffcq13txrate),
.ch3_bufgtce(iffcq13bufgtce),
.ch3_gtrsvd(iffcq13pinrsrvd),
.ch3_pcierstb(iffcq13perstb),
.ch3_rxctrl0(iffcq13rxctrl0),
.ch3_rxctrl1(iffcq13rxctrl1),
.ch3_rxctrl2(iffcq13rxctrl2),
.ch3_rxctrl3(iffcq13rxctrl3),
.ch3_rxlpmen(iffcq13rxlpmen),
.ch3_rxpkdet(q1_ch3_rxpkdet),
.ch3_rxqpien(iffcq13rxqpien),
.ch3_rxslide(iffcq13rxslide),
.ch3_rxvalid(iffcq13rxvalid),
.ch3_tstclk0(iffcq13tstclk0),
.ch3_tstclk1(iffcq13tstclk1),
.ch3_txctrl0(iffcq13txctrl0),
.ch3_txctrl1(iffcq13txctrl1),
.ch3_txctrl2(iffcq13txctrl2),
.ch3_txpippmen(iffcq13enppm),
.ch3_txswing(iffcq13txswing),
.ch3_rxpd(iffcq13rxpowerdown),
.ch3_txpd(iffcq13txpowerdown),
.ch3_bufgtdiv(iffcq13bufgtdiv),
.ch3_bufgtrst(iffcq13bufgtrst),
.ch3_iloreset(iffcq13iloreset),
.ch3_loopback(iffcq13loopback),
.ch3_phyready(iffcq13phyready),
.ch3_rxcdrhold(iffcq13cdrhold),
.ch3_rxcdrlock(iffcq13cdrlock),
.ch3_rxheader(iffcq13rxheader),
.ch3_rxlatclk(iffcq13rxlatclk),
.ch3_rxoutclk(q1_ch3_rxoutclk),
.ch3_rxstatus(iffcq13rxstatus),
.ch3_rxusrclk(iffcq13rxusrclk),
.ch3_txcomsas(iffcq13txcomsas),
.ch3_txdeemph(iffcq13txdeemph),
.ch3_txheader(iffcq13txheader),
.ch3_txlatclk(iffcq13txlatclk),
.ch3_txmargin(iffcq13txmargin),
.ch3_txoutclk(q1_ch3_txoutclk),
.ch3_txusrclk(iffcq13txusrclk),
.ch3_dfehold(iffcq13aptexthold),
.ch3_rxuserrdy(iffcq13rxusrrdy),
.ch3_txuserrdy(iffcq13txusrrdy),
.ch3_cdrfreqos(iffcq13cdrfreqos),
.ch3_cdrstepsq(iffcq13cdrstepsq),
.ch3_cdrstepsx(iffcq13cdrstepsx),
.ch3_dfeovrd(iffcq13aptoverwren),
.ch3_dmonitorclk(iffcq13dmonclk),
.ch3_dmonitorout(iffcq13dmonout),
.ch3_gtrxreset(iffcq13gtrxreset),
.ch3_gttxreset(iffcq13gttxreset),
.ch3_pcsrsvdin(iffcq13pcsrsvdin),
.ch3_phystatus(iffcq13phystatus),
.ch3_rxchbondi(iffcq13rxchbondi),
.ch3_rxchbondo(iffcq13rxchbondo),
.ch3_rxprbserr(iffcq13rxprbserr),
.ch3_rxprbssel(iffcq13rxprbssel),
.ch3_rxqpisenn(iffcq13rxqpisenn),
.ch3_rxqpisenp(iffcq13rxqpisenp),
.ch3_txcominit(iffcq13txcominit),
.ch3_txcomwake(iffcq13txcomwake),
.ch3_txdccdone(iffcq13txdccdone),
.ch3_txdiffctrl(iffcq13txdrvamp),
.ch3_txinhibit(iffcq13txinhibit),
.ch3_txpisopd(iffcq13txserpwrdn),
.ch3_txprbssel(iffcq13txprbssel),
.ch3_txqpisenn(iffcq13txqpisenn),
.ch3_txqpisenp(iffcq13txqpisenp),
.ch3_clkrsvd0(iffcq13ckpinrsrvd0),
.ch3_clkrsvd1(iffcq13ckpinrsrvd1),
.ch3_pinrsvdas(iffcq13pinrsrvdas),
.ch3_rxcdrovrden(iffcq13cdrovren),
.ch3_rxosintdone(iffcq13cfokdone),
.ch3_txprecursor(iffcq13txemppre),
.ch3_cdrstepdir(iffcq13cdrstepdir),
.ch3_pcsrsvdout(iffcq13pcsrsvdout),
.ch3_refdebugout(iffcq13refclkpma),
.ch3_rxcdrreset(iffcq13cdrphreset),
.ch3_rxcommadet(iffcq13rxcommadet),
.ch3_rxcomsasdet(iffcq13comsasdet),
.ch3_rxelecidle(iffcq13rxelecidle),
.ch3_rxoobreset(iffcq13rxoobreset),
.ch3_rxpolarity(iffcq13rxpolarity),
.ch3_rxsliderdy(iffcq13rxsliderdy),
.ch3_rxslipdone(iffcq13rxslipdone),
.ch3_rxsyncdone(iffcq13rxsyncdone),
.ch3_txelecidle(iffcq13txelecidle),
.ch3_txpolarity(iffcq13txpolarity),
.ch3_txpostcursor(iffcq13txemppos),
.ch3_txsequence(iffcq13txsequence),
.ch3_txsyncdone(iffcq13txsyncdone),
.ch3_cdrbmcdrreq(iffcq13cdrbmcdreq),
.ch3_rxclkcorcnt(iffcq13rxckcorcnt),
.ch3_txmaincursor(iffcq13txempmain),
.ch3_bufgtcemask(iffcq13bufgtcemask),
.ch3_cdrincpctrl(iffcq13cdrincpctrl),
.ch3_rxbufstatus(iffcq13rxbufstatus),
.ch3_rxcdrphdone(iffcq13rxcdrphdone),
.ch3_rxcominitdet(iffcq13cominitdet),
.ch3_rxcomwakedet(iffcq13comwakedet),
.ch3_rxdapireset(iffcq13rxdapireset),
.ch3_rxdatavalid(iffcq13rxdatavalid),
.ch3_rxresetdone(iffcq13rxresetdone),
.ch3_rxresetmode(iffcq13rxresetmode),
.ch3_rxsyncallin(iffcq13rxsyncallin),
.ch3_txbufstatus(iffcq13txbufstatus),
.ch3_txcomfinish(iffcq13txcomfinish),
.ch3_txdapireset(iffcq13txdapireset),
.ch3_txoneszeros(iffcq13txoneszeros),
.ch3_txqpibiasen(iffcq13txqpibiasen),
.ch3_txqpiweakpu(iffcq13txqpiweakpu),
.ch3_txresetdone(iffcq13txresetdone),
.ch3_txresetmode(iffcq13txresetmode),
.ch3_txsyncallin(iffcq13txsyncallin),
.ch3_rxphdlypd(iffcq13rxphasealignpd),
.ch3_txphdlypd(iffcq13txphasealignpd),
.ch3_bufgtrstmask(iffcq13bufgtrstmask),
.ch3_eyescanreset(iffcq13eyescanreset),
.ch3_hsdppcsreset(iffcq13hsdppcsreset),
.ch3_iloresetdone(iffcq13iloresetdone),
.ch3_iloresetmask(iffcq13iloresetmask),
.ch3_rxdebugpcsout(iffcq13rxoutpcsclk),
.ch3_rxeqtraining(iffcq13rxeqtraining),
.ch3_rxphdlyreset(iffcq13rxphdlyreset),
.ch3_rxprbslocked(iffcq13rxprbslocked),
.ch3_rxstartofseq(iffcq13rxstartofseq),
.ch3_txdebugpcsout(iffcq13txoutpcsclk),
.ch3_txphdlyreset(iffcq13txphdlyreset),
.ch3_rxmstreset(iffctrlq1mstrxreset[3]),
.ch3_txmstreset(iffctrlq1msttxreset[3]),
.ch3_dmonfiforeset(iffcq13dmonfiforeset),
.ch3_rx10gstat(iffcq13rxethernetstatout),
.ch3_rxbyterealign(q1_ch3_rxbyterealign),
.ch3_rxchanbondseq(iffcq13rxchanbondseq),
.ch3_rxchanrealign(iffcq13rxchanrealign),
.ch3_rxgearboxslip(iffcq13rxgearboxslip),
.ch3_rxheadervalid(iffcq13rxheadervalid),
.ch3_rxmldchainreq(iffcq13rxmldchainreq),
.ch3_rxtermination(iffcq13rxtermination),
.ch3_txmldchainreq(iffcq13txmldchainreq),
.ch3_txpippmstepsize(iffcq13stepsizeppm),
.ch3_txswingoutlow(iffcq13txswingoutlow),
.ch3_rxphalignerr(iffcq13rxphasealignerr),
.ch3_rxphalignreq(iffcq13rxphasealignreq),
.ch3_txphalignerr(iffcq13txphasealignerr),
.ch3_txphalignreq(iffcq13txphasealignreq),
.ch3_txphdlytstclk(iffcq13tcoclkfsmfrout),
.ch3_dmonitoroutclk(q1_ch3_dmonitoroutclk),
.ch3_eyescantrigger(iffcq13eyescantrigger),
.ch3_resetexception(iffcq13resetexception),
.ch3_rxchanisaligned(iffcq13rxchisaligned),
.ch3_rxdlyalignerr(iffcq13rxdelayalignerr),
.ch3_rxdlyalignreq(iffcq13rxdelayalignreq),
.ch3_rxmldchaindone(iffcq13rxmldchaindone),
.ch3_rxpcsresetmask(iffcq13rxpcsresetmask),
.ch3_rxpmaresetdone(iffcq13rxpmaresetdone),
.ch3_rxpmaresetmask(iffcq13rxpmaresetmask),
.ch3_rxprbscntreset(iffcq13rxprbscntreset),
.ch3_rxprogdivreset(iffcq13rxprogdivreset),
.ch3_txdetectrx(iffcq13txdetectrxloopback),
.ch3_txdlyalignerr(iffcq13txdelayalignerr),
.ch3_txdlyalignreq(iffcq13txdelayalignreq),
.ch3_txmldchaindone(iffcq13txmldchaindone),
.ch3_txpcsresetmask(iffcq13txpcsresetmask),
.ch3_txpicodereset(iffcq13txtxpicodereset),
.ch3_txpmaresetdone(iffcq13txpmaresetdone),
.ch3_txpmaresetmask(iffcq13txpmaresetmask),
.ch3_txprbsforceerr(iffcq13txprbsforceerr),
.ch3_txprogdivreset(iffcq13txprogdivreset),
.ch3_txswingouthigh(iffcq13txswingouthigh),
.ch3_rxphaligndone(iffcq13rxphasealigndone),
.ch3_txphaligndone(iffcq13txphasealigndone),
.ch3_rxbyteisaligned(iffcq13rxbyteisaligned),
.ch3_rxdapicodereset(iffcq13rxdapicodereset),
.ch3_rxdapiresetdone(iffcq13rxdapiresetdone),
.ch3_rxdapiresetmask(iffcq13rxdapiresetmask),
.ch3_rxfinealigndone(iffcq13rxfinealigndone),
.ch3_rxphshift180(iffcq13rxphaseshift180req),
.ch3_txdapicodereset(iffcq13txdapicodereset),
.ch3_txdapiresetdone(iffcq13txdapiresetdone),
.ch3_txdapiresetmask(iffcq13txdapiresetmask),
.ch3_txphalignoutrsvd(iffcq13txchicooutrsvd),
.ch3_txphshift180(iffcq13txphaseshift180req),
.ch3_txpicodeovrden(iffcq13txtxpicodeovrden),
.ch3_rxphsetinitreq(iffcq13rxphasesetinitreq),
.ch3_txphsetinitreq(iffcq13txphasesetinitreq),
.ch3_eyescandataerror(iffcq13eyescandataerror),
.ch3_rxdapicodeovrden(iffcq13rxdapicodeovrden),
.ch3_rxmlfinealignreq(iffcq13rxmlfinealignreq),
.ch3_txdapicodeovrden(iffcq13txdapicodeovrden),
.ch3_rxmstresetdone(iffctrlq1mstrxresetdone[3]),
.ch3_rxphsetinitdone(iffcq13rxphasesetinitdone),
.ch3_txmstresetdone(iffctrlq1msttxresetdone[3]),
.ch3_txphsetinitdone(iffcq13txphasesetinitdone),
.ch3_rxdlyalignprog(iffcq13rxdelayalignprogress),
.ch3_rxphalignresetmask(iffcq13rxchicoresetmask),
.ch3_txdlyalignprog(iffcq13txdelayalignprogress),
.ch3_txpausedelayalign(iffcq13txpausedelayalign),
.ch3_txphalignresetmask(iffcq13txchicoresetmask),
.ch3_xpipe5_pipeline_en(iffcq13xpipe5pipelineen),
.ch3_phyesmadaptsave(iffcq13phyesmadaptationsave),
.ch3_rxphshift180done(iffcq13rxphaseshift180done),
.ch3_tx10gstat(iffcq13txethernetstattxlocalfault),
.ch3_txphshift180done(iffcq13txphaseshift180done),
.ch3_rxprogdivresetdone(iffcq13rxprogdivresetdone),
.ch3_rxsimplexphystatus(iffcq13rxsimplexphystatus),
.ch3_txprogdivresetdone(iffcq13txprogdivresetdone),
.ch3_txsimplexphystatus(iffcq13txsimplexphystatus),
.ch3_rxphdlyresetdone(iffcq13rxphasedelayresetdone),
.ch3_txphdlyresetdone(iffcq13txphasedelayresetdone),

.ctrlrsvdin(iffctrlq1gtrsvdin),
.ctrlrsvdout(iffctrlq1gtrsvdout),
.coestatusdebug(iffctrlq1coeregrst),
.correcterr(iffctrlq1correctableerr),

.debugtraceclk(iffctrlq1debugtraceclk),
.debugtracetdata(iffctrlq1debugtracetdata),
.debugtraceready(iffctrlq1debugtracetready),
.debugtracetvalid(iffctrlq1debugtracetvalid),

.gpi(iffctrlq1ubgpi),
.gpo(iffctrlq1ubgpo),
.gtpowergood(iffctrlq1gtpowergood),

.hsclk0_rpllpd(iffhsq10rpllpwrdn),
.hsclk0_lcpllpd(iffhsq10lcpllpwrdn),
.hsclk0_rpllfbdiv(iffhsq10rpllfbdiv),
.hsclk0_rpllreset(iffhsq10rpllreset),
.hsclk0_lcpllfbdiv(iffhsq10lcpllfbdiv),
.hsclk0_lcpllreset(iffhsq10lcpllreset),
.hsclk0_rplllock(iffhsq10rpllfreqlock),
.hsclk0_lcplllock(iffhsq10lcpllfreqlock),
.hsclk0_rpllsdmdata(iffhsq10rpllsdmdata),
.hsclk0_rpllfbclklost(iffhsq10rpllfbloss),
.hsclk0_lcpllsdmdata(iffhsq10lcpllsdmdata),
.hsclk0_rxrecclkout0(iffhsq10rxrecclkout0),
.hsclk0_rxrecclkout1(iffhsq10rxrecclkout1),
.hsclk0_lcpllfbclklost(iffhsq10lcpllfbloss),
.hsclk0_rpllrefclklost(iffhsq10rpllrefloss),
.hsclk0_rpllrefclksel(iffhsq10rpllrefseldyn),
.hsclk0_rpllresetmask(iffhsq10rpllresetmask),
.hsclk0_rpllsdmtoggle(iffhsq10rpllsdmtoggle),
.hsclk0_lcpllrefclklost(iffhsq10lcpllrefloss),
.hsclk0_lcpllrefclksel(iffhsq10lcpllrefseldyn),
.hsclk0_lcpllresetmask(iffhsq10lcpllresetmask),
.hsclk0_lcpllsdmtoggle(iffhsq10lcpllsdmtoggle),
.hsclk0_rpllrefclkmonitor(iffhsq10mgtrpllrefclkfa),
.hsclk0_lcpllrefclkmonitor(iffhsq10mgtlcpllrefclkfa),
.hsclk0_rpllresetbypassmode(iffhsq10rpllresetbypassmode),
.hsclk0_lcpllresetbypassmode(iffhsq10lcpllresetbypassmode),

.hsclk1_rpllpd(iffhsq11rpllpwrdn),
.hsclk1_lcpllpd(iffhsq11lcpllpwrdn),
.hsclk1_rpllfbdiv(iffhsq11rpllfbdiv),
.hsclk1_rpllreset(iffhsq11rpllreset),
.hsclk1_lcpllfbdiv(iffhsq11lcpllfbdiv),
.hsclk1_lcpllreset(iffhsq11lcpllreset),
.hsclk1_rplllock(iffhsq11rpllfreqlock),
.hsclk1_lcplllock(iffhsq11lcpllfreqlock),
.hsclk1_rpllsdmdata(iffhsq11rpllsdmdata),
.hsclk1_rpllfbclklost(iffhsq11rpllfbloss),
.hsclk1_lcpllsdmdata(iffhsq11lcpllsdmdata),
.hsclk1_rxrecclkout0(iffhsq11rxrecclkout0),
.hsclk1_rxrecclkout1(iffhsq11rxrecclkout1),
.hsclk1_lcpllfbclklost(iffhsq11lcpllfbloss),
.hsclk1_rpllrefclklost(iffhsq11rpllrefloss),
.hsclk1_rpllrefclksel(iffhsq11rpllrefseldyn),
.hsclk1_rpllresetmask(iffhsq11rpllresetmask),
.hsclk1_rpllsdmtoggle(iffhsq11rpllsdmtoggle),
.hsclk1_lcpllrefclklost(iffhsq11lcpllrefloss),
.hsclk1_lcpllrefclksel(iffhsq11lcpllrefseldyn),
.hsclk1_lcpllresetmask(iffhsq11lcpllresetmask),
.hsclk1_lcpllsdmtoggle(iffhsq11lcpllsdmtoggle),
.hsclk1_rpllrefclkmonitor(iffhsq11mgtrpllrefclkfa),
.hsclk1_lcpllrefclkmonitor(iffhsq11mgtlcpllrefclkfa),
.hsclk1_rpllresetbypassmode(iffhsq11rpllresetbypassmode),
.hsclk1_lcpllresetbypassmode(iffhsq11lcpllresetbypassmode),

.m0_axis_tdata(iffctrlq1m0axistdata),
.m0_axis_tlast(iffctrlq1m0axistlast),
.m1_axis_tdata(iffctrlq1m1axistdata),
.m1_axis_tlast(iffctrlq1m1axistlast),
.m2_axis_tdata(iffctrlq1m2axistdata),
.m2_axis_tlast(iffctrlq1m2axistlast),
.s0_axis_tdata(iffctrlq1s0axistdata),
.s0_axis_tlast(iffctrlq1s0axistlast),
.s1_axis_tdata(iffctrlq1s1axistdata),
.s1_axis_tlast(iffctrlq1s1axistlast),
.s2_axis_tdata(iffctrlq1s2axistdata),
.s2_axis_tlast(iffctrlq1s2axistlast),
.m0_axis_tready(iffctrlq1m0axistready),
.m0_axis_tvalid(iffctrlq1m0axistvalid),
.m1_axis_tready(iffctrlq1m1axistready),
.m1_axis_tvalid(iffctrlq1m1axistvalid),
.m2_axis_tready(iffctrlq1m2axistready),
.m2_axis_tvalid(iffctrlq1m2axistvalid),
.s0_axis_tready(iffctrlq1s0axistready),
.s0_axis_tvalid(iffctrlq1s0axistvalid),
.s1_axis_tready(iffctrlq1s1axistready),
.s1_axis_tvalid(iffctrlq1s1axistvalid),
.s2_axis_tready(iffctrlq1s2axistready),
.s2_axis_tvalid(iffctrlq1s2axistvalid),

.rcalenb(iffctrlq1rcalenb),
.pcieltssm(iffctrlq1pcieltssmstate),
.uncorrecterr(iffctrlq1uncorrectableerr),
.pcielinkreachtarget(iffctrlq1pcielinkreachtarget),

.refclk0_clktestsigint(),
.refclk1_clktestsigint(),
.refclk0_gtrefclkpd(iffrckq10refclkpd),
.refclk1_gtrefclkpd(iffrckq11refclkpd),
.refclk0_clktestsig(iffrckq10hrowtestck),
.refclk1_clktestsig(iffrckq11hrowtestck),
.refclk0_gtrefclkpdint(gt1_refclk0_pdint),
.refclk1_gtrefclkpdint(gt1_refclk1_pdint),

.rxmarginclk(iffctrlq1rxmarginclk),
.rxmarginreqack(iffctrlq1rxmarginreqack),
.rxmarginreqcmd(iffctrlq1rxmarginreqcmd),
.rxmarginreqreq(iffctrlq1rxmarginreqreq),
.rxmarginresack(iffctrlq1rxmarginresack),
.rxmarginrescmd(iffctrlq1rxmarginrescmd),
.rxmarginresreq(iffctrlq1rxmarginresreq),
.rxmarginrespayld(iffctrlq1rxmarginrespayld),
.rxmarginreqpayld(iffctrlq1rxmarginreqpayload),
.rxmarginreqlanenum(iffctrlq1rxmarginreqlanenum),
.rxmarginreslanenum(iffctrlq1rxmarginreslanenum),

.trigin0(iffctrlq1trigin0),
.trigout0(iffctrlq1trigout0),
.trigackin0(iffctrlq1trigackin0),
.trigackout0(iffctrlq1trigackout0),

.ubintr(iffctrlq1ubintr),
.ubmbrst(iffctrlq1ubmbrst),
.ubenable(iffctrlq1ubenable),
.ubrxuart(iffctrlq1ubrxuart),
.ubtxuart(iffctrlq1ubtxuart),
.ubiolmbrst(iffctrlq1ubiolmbrst),
.ubinterrupt(iffctrlq1ubinterrupt),

.rxpisouthout(rxpisouthin_to_rxpsouthout_q1),
.txpisouthout(txpisouthin_to_txpsouthout_q1),
.pipenorthin(pipenorthoutq0_to_pipenorthinq1),
.pipenorthout(pipenorthoutq1_to_pipenorthinq2),
.rxpisouthin(rxpisouthin_q1_to_rxpsouthout_q2),
.txpisouthin(txpisouthin_q1_to_txpsouthout_q2),
.pipesouthin(pipesouthin_q1_to_pipesouthout_q2),
.rxpinorthin(rxpinorthout_q0_to_rxpinorthin_q1),
.txpinorthin(txpinorthout_q0_to_txpinorthin_q1),
.pipesouthout(pipesouthin_q0_to_pipesouthout_q1),
.rxpinorthout(rxpinorthout_q1_to_rxpinorthin_q2),
.txpinorthout(txpinorthout_q1_to_txpinorthin_q2),
.resetdone_northin(resetdone_northout_q0_to_resetdone_northin_q1),
.resetdone_southin(resetdone_southin_q1_to_resetdone_southout_q2),
.resetdone_northout(resetdone_northout_q1_to_resetdone_northin_q2),
.resetdone_southout(resetdone_southin_q0_to_resetdone_southout_q1),

.rxn(gt1_serial_rxn),
.rxp(gt1_serial_rxp),
.txn(gt1_serial_txn),
.txp(gt1_serial_txp)
