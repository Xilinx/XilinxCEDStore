
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2023.2"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
grFagMniYm1tGWTRjQXFHLc/TyirnHUCzhk5hRPvg8qDIZ7zqCfDjr4HtQ/0FDfqIt97QEy1G2NF
9/t9SD5NgnT2cJ33Myl8XcN9ALej/6hOLRJziSvpXQcmzGAS14T9cyfMYf8mTlneL2MZov86IFWM
wHzMz8as4w3LT2kA1tr9z5Q9WiYVc+Xgl33gdk2bFgW0iMppigXbdKTK/ipo4WFtTu5uifFBZD8Y
MUaDGqs1eaD/qeU6XQVLBuBRbmtW0HbCP57hoSuBEUUK1vylVNYnmJ+TGp/fmFiCEHP8sEp1VVar
1eeXCSMRIg9UpzWnRUu4BUObFppt6ZeAxewi7A==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
sPJDQN5PzCow3WMEDHilgqdRL5MnqiaZhhG209q6Q+mDo0Wj639OXcAcvl6T0Qr4lamYnNLFYxNL
QcLZOyoxxhzoFqO8hz1C6cTqrmYvGWcNDhRj6uGee9tMAM4VAbO8UjlIF9XlycQHvY0MZJ7i3log
7RleJQ8VyQCdd9KwTQZhh/It7oRLEGGQNGBV61M4linMob99xBy89YO3/1STlE37AgFHCxxvIV1m
AUomaaK+bVOV6Te5glPDHX0YM8ohdltnByUO6iFQ+Uzl12jvtCZqBP0R+zxR8XCgA1/TKLXcJav/
Ax0Oo1xzVErjKZbQEDkJtnNNo79GcODwu8SUyQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
d1WZiNNPMj1nVeKx7u3y3fR7rJrtjMbRwrAeEb7kmcLXWKDEGN2h0M/K/QoK22+FyDFJFWrp31Ya
uq2Gn+sCRoaSxJdySdjue1xptoUNrmTvNhBKWE6crNASQ03vj7jyjDcGbsnqusFyRM8mxXGbBmfb
0b3OLTaUxapwIzix2io=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
oN6NzCQWYpX8CBZiwOKQRrkD8MvicTzgBEmOVZiF3b68Rkp/UA1lMrgIBxAsGNsGyfczvGwjrfGg
/YOm3SPyR6B4ADGtSEZUDIBYEv48SX1XXiME26F+FMiVJ6n+AYAjaB4s/3/H8MH+XAOQF32+hROh
rS4Fuw4vJY2OacS2JfTJrVO7BXMVRNOgYRiT/mHX5NrY1TCZiPIIcJX8mbnuvT2Q/Qo/iu5Gwlu3
8obvpmTMd6Hc0FSCiNg76iOeZKQhtrepaxr/X0N/jAfuAZT74ARxSWWHI7iuFCQ8yaWcL0ut+DEt
BQbmbvLFP9uFXkDFUxJVB0g+tES+BvE4omYpAO7L+Ot15sY4j4P+2NEmZKUVAUNrhpVI/NO6KAdF
LdJ7+YOmpEeu4dcxj7y2VbLzJimWUWW8V5PAk2bvHm6n97vMEGYQec86+N0MCkrs5UU3IF4bnoDz
FMYcowOG4jTG9nfDhia4DEaJXhscICdNDQotl5qmTvq+zGouC+p//HIA6wK2ZJ8KitTSSnG9L/nC
IWaB0q9EH9AKiAQIlZlS7Ac9hV4JJbcNpYTuAd9c33DdbiE/biO8T2L2qCkbLqeOqouXSugUNKRo
a+Jn+1GbGNznhantydgBJlWjTGAWkPg5gTx+KnBZgAu6OOpHyL2aywR/Xx0T2GKiQ+dorWdLLULr
dvVVEWAUlb+DlzCbw8Y63HZWFr1cLCKqgWFdPxfGff10OPjg0lZvU2YDIn4lYCMprGtyZl/IQe5G
MXxd1c5qtuaej9Fxc3x50CNZQyp2vdGLGi3rvfoEtC80sqt0gR2dW6D7cW9V8gzGATN7LLfUA17x
OVDyV0zQWzpqDRGIAV/aLZKHfi9Q3XN2rFLFXmygNdu9+xKC6622LYGZitMyupOTDFgqNhi5OiSa
ETgZ866aDrMuAyGl5qRxA6Q7hu8+pIUdySinZt5/81CGHr/lP/h6St6qITWcNDClLpjks/PueZ3v
LMv+gbQXpiwbNvZ2f+RLTvTc68JT/7U5a9a8rCpowN5czdDCKcyp5EXAYZ05IIaOhEan0CVcj5Bs
kf3P2BYc/NI1f9Ac4LFiV2SskpJo8YrPWrMwRtKEJqeJZtAraYWPqR6ZDPYyuotLnxPSntuHYSxL
DVguuet1D+2Dc5cj+PsRYuzHEKwY/lStVsFb9UyxtMWMu1fb8duDVZr9EaB7qA7bcC2OkaPgqa00
LbSWlLfrp1o0/aScTxDC2Qz6LMW4HVtEcOROAzrFo3WFjbhqaXKLht9XT9XsoB132oXEFdufhVvr
RW8kCYbjdjUuu2go8wo7UkjOWhliuESR9LS6fM1phMv8eMdvTWIqXeBK3aLKgUL0vZs9MYKh7Anq
OLK7g/2Xq2njTA4LtBifk7SbYiPFNWUlGp7gp7+9iOzk3FcQFcr4sq/DVc5hrjMp0+c+BJlaCCdl
nPYbIoQW3IWY4Md7m98kyAswA0kmRDtd4Jpvw8wnwwk3opDE6Fw9LvMXIjVHcKOUs9JttVdZNgtg
3Eq5ex/en/Q25bQj72xDnxKN3dB3GeuJMQnEuPj/aHPXvARPGy3nY47JuXYqT6eBgF6vys+XjEG1
A/C0rZPhN1q6SG3j4YKBpIQAHkGc8h3AP1GjMc1tRqiC4i2+KzO4g6mlp+pK+HW9bpQzVZB8eYgG
6O5U2RGFhj9VwU4U3KTcwNopVBWmbuPclJiZtXvYSidpfAycjPVk8xZ2jw3KynglXDg7ZyoDWyc/
EYY93vaUnRG520n41pU+J30j8dbVFv96So9qIEwyHqa+4toLQ2vJCjI7ELCEnPpivBuDe/Ok55tF
ZOCaoBvab5/VPPvJyDLqbbKpQJLzwRCs+0tZcEmFARa8QASnXIm3LP55LkNKLGIGHLlj4jVLBj43
DzSxPiru1oEn+oqzFadfDN2sFxAcMNLAEioF9/g6gQT6V+6nf76/HfhMQ9gKayWP2w4nlxzUGBK6
RAOlGXsOgUdB0g4zE45TbLdzLp5eAJDaocnZEmUlKkWwYziSGfKQWbPhPDa5smKxkjgW/FQbDt9U
duKRwTp76D+JIpZ9x3E2m5vTxznrS5Vl8P1Ebm1ItDV7hntoRfSUusDpvaTdelcazC8WA4Uzh94N
NTXEXec/BD9QS8if2GvVTfwGrj4vNo/rIIhM2ZSqlekCtF2f5yvCrL2bB0ysaM+Urnh/T4F0gp3A
tLQqz8okeuTc6cVMV8BUvJMdzqjnx5mI7jN+BAY/8Juo6ZL5DmaRWFgxuZOF86mCxnnM0v4N+7+C
SRC2iB07zuvMKRTS6lWsKdWGH1dLPa0WuHDxhWWcAqZ0iDwb8lF5QqrCxMd7blTjwMzTEQz0Jej8
nhFrqf1mBZcId9qydVxWiSu2lXiRD8QTrcXKTWCVXzppHIqUKOtkRNxf11MLfkrCqOl7RB+D8S+O
+5O/Mh+cVzMrVtehgBqs7rre+wrzMtRCiAcqoj7LxA1k0+Z9M6CnikczkaSR46sdkmEZHXsWF1Ny
IMdE5WWOZFMtITEDxiE7KlJBAoPYxC8UT/epf8wcyrZ9AqXiOyH4xADfuq+59mcB4z+EL8ZCrKGS
TT8DXoL3yM8FYVhIQ+9Pbnm3aFxkwcHXjxGTx5fHMF5Lk/IW27G8HsSSPuib7a6l4QLcFz2fvGZ3
ntfq3nh7x2Z3kHbAJe7+Og0N55BA/Nx30JlW+YBBB7YiWyJ0jkJL4BsHJyF8pWfHe4i5ELUy2ScG
xSHbzUHPuO6MypPMLRANBtmxYa/iCm8CI3aqba1ujL/H0FpvyQXXeEgynYKmrACofxc6Iy7lnfE2
f2jsY5F3t06zViLOIh8449t2haQaFen2JTrtFVb5SpHy31uA5Lk3s8LC9xoZzZJCCrE8BAEKb4x5
V2shXl++QszR/Pr8wjtSp8SoTAxFtUwhN5SXFcTE1SpB899mDfSwhkSLzAagNMRuudaJR6YeN1HT
njJHM2jdnmJ3u+NCgtbY9HgwDUBSQqZ4sUvhlsuUN2xlmYX4sL4wC7qBo8Eckbp0u88RQ+0Tc+1a
mTGPbpY9prRwtAyCRuKV5VbyLHIcg3mw85inyGLOAvuHp6I6ek6J6hiEZBWJKJmzyANnERZFIdSz
Gphx/HJ2ZLaSAByvzH12nkyw+vFFL8aMdE3QczWIHFY0A47rbYmisLKkhryFzLfHnCnD5McMzyey
Rg0LvUhvm5mvau/IdCllojY8oUwhbzedgqp8pQuqFNC6ofVEHCKGJ5F9kK0rZevaglojbE684/Xp
OX7KQJnfsDzcEbzjEOmHfVXrd91RGbkeeeNh0djqVEbE0LyzNvsu0EqQvpwnSj9RRAbHfBE++Dsa
GkvgrX3f+DxfDN+XlVrkflUW3ySxj872lGPw+fLz1L+6EODESZMGnRp26avYLTPKu0YHDxihx63p
reghV784xPJhP5lboNBuEfyNwmQE1VK9+AhxfDAHpiDY0nRzN80GYiSw72HOEodnLYX4RV9KbBy8
oQi0g/5tjCiSjRlWNw076JWgf3R1CM2g0HKTLPPbGvr+DDdVLe8lXK4F+4dLk8rvLK95+DZIvLxV
ryD4CBOu7PMWrf1J6ekLysWIy8sKeSL/UL384e9qfQnnX1qJ6jvH5UqQkpUdqWbkXU1cP8fUWsD1
dZSVlEh25Jo/bSDqRoqnFjtuwDFExIcdRoNKxshTagvGpR11ijT7zVk+FKLWoxOU3CjuBLNl1Ln6
DyXq3RHZ5znADm0A0EsFgHJkxBLdEF1SKy48kT8cDZlrCs8/ofGo7QYMGA0tj6c1+uMzlpF7XkTx
poSh7nrWqEWMlSPbFJE0qvV/+V7i+xSJL2sELRhsfxZ/ZSydiYIpHd57Kr4LH6hypQNFss2792nJ
Di0Xv6Dfg2q19rGGJVuiQshxxKSJ2Voq95a9u2svgnSV4iue+7jxvwprNrYx/SxIw5wS0/OBgnDp
XR9JayPQc8IRD0RyG1ULkeDKbZMUb7Y8wz9ukf2s1riEZ2DYSDLLV+ITHB9WoCjkzFlWSLGQHKTN
2BB7nZWLbVYeIH4MxqGZogJynjOvGJ8xR8Ll94pzDe5bbpZ0kpSqgkeFK6BegRSuBPrT0rrcn3CR
RLTZQ+Z1PCLYRAIHmswP12PSq7bpgaNPiTwn80lD/S2b12IRAArl3vsHZT2RzSi6TM7cDSZBVRyt
xf+1Taob5W1p8OiCTI9rxPn7pSSl1z+JQOgKbJ+HRn1Plv0UQWiwk5A0RO3sxsEkHPnKyopanpNv
E/M0iIru9+lYdV7R1w0FAVH+1QxUkGHJzKbV+lfwDTefVnRCM69xNJJYaWAfrF2hAN3BypAuFaRB
ni9EXRYqWvDxy/gq3xh0a0BIN0BzkBsLLhA9maN9aEJ6i93uTVvn3Uu+Ajc8u2WMrYiYKl/wGHkz
BFkRV2bEfuX4SoFhXRpjADiiNjLvEE/Mc0gw1NqQcLZBb12s0ygaNKLYivN1fcEZC8cjZb8N07Wv
xBzA3AWeB9QX6JZMzmYhkVxWGPyhP/RXHXUQ3CJC535KOIiDuLaKPDupRNLLbq0beq0BJ3xPYfFc
UsKTAJFVsTTrIjoC8XbL18taKQYq0AF4USMZhcmW23vkMQvktOBpZIt9UXJGov0M8t4k6DF1Chs1
7jrR1OKf243FOW9+v1AVY3mefzTSGK9bKNW6JRve/ci0/vbS45K0ap4SgUW0B9Gwt7KsD8xvi4MU
GerCMrSFusHX4QXllwjxmlETRQ+Czq4kQLIFL9nlfsr2UsvO6BNx1NMxath5vbX/OnpI5aGuR8Mu
V6RyMs2M95NVbH3MyxsW/W1scEjwHwHV1rTb2TM89DwGT/Pl5oHHCGRaEcZn5Qzfd1dqlos2gi7/
/Aml7HaKSd0CEot2QpzFHfos0ezaOPceS0uTFExd6kr+dWUvENrXGGZ4qhKyFKZeFcCqX5jOXmBI
CmGAR5gGw/DAo/9C8rtK9e4i3gbK8V/LvahYQZwuE1Go1/ymQnOFjTHIuJNrm+pBuSS7If2bBk3D
C5+mWE3amksv/OVN1ueqSBWpbNlswHfymIEY0JrHhHTjJwGk7ksUf0x6YNdXVIOGn77I0pNsFmsf
qadrhdcwMaBQmUMA4t7dr5iFfRUk6bppPWmwnhfjaBFh0Ceis/ahCRQaFADdtKjcZryq24AepB1Z
V4RoNVWqWg8ZmrbHSHNJCI5X9eMhHQlo1I4lZful5jpyOF7vc/GwUlJRrlZ8mKxI2z3feCQuTfT+
wvrfFMkUe2u3y3Nzq6Sl2cuuSVrW8Licq/rkAQW5RYzmAF8AOj5xgZ8/0G5TNvea1W651jVNxH2g
YkyYkUYeaWN0ljUIHhGctCi0XtVuIQDC16GXFV+fW2DFAp0+DaupZnh0YoPSx8MLbOXpu+FnuOLy
awYQlCym3FJO0YQteiVgJ22IzHj+3SVSPj0TZiY2HWBvlFRjXLj8i+pS/Nz4eCnVHfdxmZyVPFE+
/THjpn/zso9Z6MGUwCQUXLnlpz/09LSQWZdWMU9NnwW12jQBDdtKSzZHGvnF9RZgwmiuMUMrMURx
ALVfKyPUSlNoKnClBFPwTQPL51ViI99/wDfqRzhpZo4TchTCHd2u5kQNsbEu92/bI+McgCa7KT0Q
GrkupNlpnwJDiafIRyspRETHk+Rlkrz/SqZ563V+SzrSiMjHf+RnMfqcnxlnMfNBlPYuN2tiNtdo
kwMqKcXqf44YyZuTXsVMbXWA8Qf/X1Ehtba3Za7iVHkkt8Na9/YJ2GqYa+SbRcZcofY+99TBssfn
wVNSri+22Ogt0Aang+m4Jyc8B+j/3IeX1V7n7XWQUXiFdRlISHsS+1o4X55AfmzKGO93on7AnJfG
aWvhJYinUGqprmlJEbQAFXeSBquGOQtHOxug/uIyc4A6yiiV7c5nnEmU06K6BZ9+d3gJTw3M7mnD
27szsg1nPT1eJgH5Hj6iieMBV9s9B6ZMtFujv7U0MdDI2ycTkujrQ691sOcGaUT7d3ty/ZcCA9Ff
V0dhYjXVsb3SNn9/a+rIJfIb3C+c225B+QFpoJkb2nYuo57baAM/gECUS2W8cWxDeCvlEQYrXPEz
1aPcX1rfAMnPjWVNW33elC7Zy1pkBVRlTkyaYteR+BV9S3jXR4NlQDw4UKGZpsP7exTObycSckV0
SMqB+6w8t9fRke2KWLImohqyoYpSFZjSydjv8e7CBbRMLY3zBNV9mcMZPrirj8ZTFb5ZwjLY6YC3
5XF8PTxReLg0VQslS7QDuS4CCbHcJFc6SA5lcDBF+FX6E20Ubdum5zPAJAciOmS/Mk35LnsBbsvM
6vcMFEoRimDPgPqBv5mVU7gBxEMBVTSV8nL8t65uxwZXzfTURTSpqo6Dl7oFbuOXC/Bj23dqnek5
AE95PovwzVe0Gk+k2z9YWuqZWw2FSNth9l+KmTw2hazXEW54ebvxiGoPrRZh+vs2cs04ZFQdptfK
axb2IWxSglNvZbz0Vc8Zpap0RO0G7+C24It1ZJu5gPp1CTLGF/69Yp7/FEXtcJWJu3IY7T7hQ+n7
0klxYfkqTQNQAdLRJwPyxWb6dF9/7nby0keXS0YJtr55BwCBXH2kn4HPdi0ehlKg4qK9KH2wBFj/
EdBYQNvEqCAI1awwNSg41qurtkKH/d/85DHBKTjZ5XsLzYGg/FUud6gTUNMlGI8ffAiS04nwIza3
1/vM0lr2+2IOci7QQLkb2sTGe9ldyYka5iZ6UJDs3Ja56xmH1wMlPdHNnmsQRGrH66qMUQVAbxPO
heSwNegVcFQ5xbEUcCt8mamBo1iv2xZ1jA1v8u61eF5DjZGKWzDGwIp6eL3ZExecXkvklpZkm7b0
vG0bVXM01id/QaMPXmXEltdn1dDdXTj5ekAer3efJ3T/npttIvZX6Z8NfP+jmlKCuQOsnAogZbzS
6jMv6FtdXEIObJclQlcPT5NzAwpOoFJMfSCIXfddXfwE9TU12qd3mO3ZN/A23Tv7IZAiVoUY4oGh
lC7qr7d4LCps1RmN2/nQyaPgRu295jFOUV+ykz+1pazJ9UPf38ftSpZHeDiNvJLZVbsyOlntx/pq
pxpVf5lwgTU1RZzOhHIYVMqHeKyd+B3MS/72flZoJ7TsAXreryyd26rGln+aH949jXgRbEhuaLEx
sS4Pu1PZKek9jWP6gqjBQRz/lKhY/+JD/Wpfto9rZi/+3TzBZhA+Ey9TDMmZ0Vp5N9EZ7F/JVcum
aefLL5HY6ZoO3HqYHbKu66DC5vjcKj2mZJxL0p+tZIrI8DgejeG4Ccy2R0GEmXrLjBD8vQmx4M9I
gzNLDGicgw7IaOV/6l/1p2rLo5pqFYud2xiJ4xhkT5lWowKlkMGNOmPhCONWhsA2bTjZDTSD4sLQ
F+UojRfP+qq6t6cMqRVTRFvFKRVyV2t7qyU/+K6WgpkVEaeVZtoyqRzy4FbWOGNWselzDvFeVaNx
OjE+955V3PJERwuKNHgGwVKuN1UPr7Pv+bVoRUtdFrs7hkuFo5qywnnsZR5Fl8xDe/Qomu30tGZN
v42L3jACH11GseDq7aVKcUG7UtoEPBeml80WlNjzecOgB9O9o9mHIdGMs6+uRk/VNCgb6fcZyRAw
hpG6TeqivNsLuJuH7Ux1dO2Tb/Ku4eHB0QzBIRFeyMkzSzt8ZXKaNxFi2/8i06hArUS5hmyJX2WW
c8jyXMpy2G/sByvb1lfchPAXlOLobk/KhGKJr15XhGLoF6ib1yNpu/AakO7FxwI2fboZCqVJl3t9
L6fi04Szt+d4EAnrm/UKAdKo7fX/j9vgPgUNsI7Nni/m7ve1bamDemBDEW/bgsEojT7Jqm4yibM/
jrwFDkBesB946rz94/UAMF6IpqMsspF8+xmwxQaT0tWb1N8QZt0rn4WMRBIo5tc2wRkpHDNUmjPk
T9PqNkZ733WLZllJSw4kzCq8QavhaJPrkPXhsguzJtMwyvBp0gd3zZP6DgWa+oqFHXD3czUavceV
V68bXgF9b5XhPC8iFy6wnsIroAUI9ULneCbkX8ypJAygRwjeziWb9xVtET6aav/Yk9jnl2bDzq97
XJbi/Hxi18x6XK0pV4Wi0qJlGcS1YutfrV4dn5Q64LP2uMPiPPO+W2tm5QTS1SFCK7KOkFpRXqUK
nfU1ps70/3CiO7ScSylO2w3m1xBzEASDpUrr6Mcg1Rlw02yCnFXrueab9C2WuuignEqAF+gNLJFB
64W+MNCIiGgXOF77GESypdOO9CLHPs+GpUuq7EONbuWPImpLXJikPhSOpmbqx37OHgwWfaWf7VQm
+FXBr6HKUSjPwadbmocO9semUSPL1pMAsPnArobBVlolkEwFoKCuJrtdC8QFTTQ9bYlp7jNvU9MV
U5/tE309WVkH6TKenreTw9GlrF9jPHRifmz4GfEl7dvQZrFg92sIhCqZFDlxrEcgvyHUJxYaN5kG
OWZQ+wutv54+jun1pWnvqD3AqtISTfdEaZw9163w/ZXbXXMz33gfLPhTTDVEFkIzEREIz7VEFyII
y71s1Xwre9S+aFlp6VJ64YF6AIQrA7QLxJOIsk7yll38m8NhbKo/1z/F4mV8HRs+C/qFFAbPFaXu
jSv3hVk1mgMEZPWwfRwOX9CrtjBD3WQ6MoOVz0oKj5gDqJUTrqFCKKKICydFSNtNWebLmS7wSjLa
28i7gsg9wxvGUtTpdaFkpoQoFS2EfJPOAM07ufH1I5eHlvAMV8FtC+H571dJvM/Fmkr6rrJRMO7w
YSNhTJ5s4j8uxmEDfdObmb1gosQ36P2KjfHDzmiqUVuipjqW/IIVq/qJS+Ec6U0G4fGdDximRga9
OTGDGLu8GQC6H+kqAm8NbOfkPXeslRGx6rcTHtaX7+chDY6hXFNx14q2AbxzjIbImdE5HZPwnfPd
G7TV/Cs3Tmv9hMRE1KsTRXeZDiLYcHMGIsrmvmjMIijPq+8L1BfkCPSpq6T8paEJMP1MueerKCMD
rhEUnJkBn6yy4NkfTK4fYDwh9c8ZzMbWvwNKptDLRSu7L9/8qc1y9Kf6PZufcgoCXX57cDjO6ApG
9ZTWEiN4yohXUODS9kY5QdNXOETpAEznGsLbZdVcfRrAV1pZKHSFDNxIHisaj9ytLcwFRd0TCrQK
fxnii1n3o4gKuxzTUcCN/RaiSUEzfrcNa6eAIkJb6Sdlfq4g+XeatlUitxiICtwvCt1pDLhXHVPz
AkMcZvMcdmAbOAGEEfCUGuAcWdGpl+CqtYQJwVGvoeRAscZXzuWgKAuMpVwsn8z2vY2duB6cfcmq
IdINZIGpBqnnlc7qGrEam86oAeAMi+3BjVzhgyk3MttnP4+vMcjGIMOO5QsRMPsdpt2aaeGS3oll
iDY7ZfvSXE+9mbiYwIVu8OjlxzriCXQVW3ljEpLThX+QhI8IMeDbgjXC/IaSS4CRcge08TuYoSHP
TeEn9z6JYW99qE2AhEtXafrlLVruf/sTxsCDKNiRcIJ+vPNIhBfJeOfXprvFO5UyF6EAtU4TJ/0d
vvkmvLGOFBMZ/kakbDRDAGG4TwLb1trSSyhPb2bA6Zo2ow8dgW14xq935G2BsdNXJKAwegpGh1mh
fqABHvYj8YcXRYXET2QvY47hNufvPDa423xmaB7HpXwDHWZDbSpJIQO25x4Fn9VqnHJ5Jng77TNm
KAwUWqoEaWPEN9fJwCktLmL5W0hywVbUEym0fj833UwRifTS8GbOHKkmZS1o/J8P0wlL88wcCoYV
9UZUWz/fVriVSQpl18ZrC1bXhBUdfyNU2x6EpgUkfEjAyk2+Ehv2z13vFbksKYbG087EOq17hVhd
+4DrYVE1mLLjHpJmiHQ9pmwLgWl87dAyPDBiBSkGiL9rlY+Fb8ky7kTyXsHzVaSDzoGp+wNyvv6m
UOJE1OlNynSrxoyOEx3fynqS6/Awy3LGOmJalP8AYhQq82SfEB8K4OW+kLEOSmf6CT3u81b3GhPm
NxaZTEsKpqzOAUCO46IydSrz24AohRh0byKJby1EjeuK14kBLeZOjDu0jbyh/soHr5OOdqzoZnM3
m3ORUWopFDeY6T/LNhc7qisAq4NG+MTezXk2IyG5eWzdHLCRYDdC1M4PoYruzFzZki+L5zqnYzVd
MxHMxi99N+C112raetxc2lpOJBUro36HAwTHpnsjQjqY/T966YyrXHDgQVJtMEqJGfTbrIOScvN+
qseSISm5ZGIDIo+Dt1ipb81roJiuDPfKz6wQfvhyZqmSSpNqbty9rr9HRYZDpqFAlGOjSB5AHmlD
vJRoW+8kkZTTK77SYoAmlZOn977ONOC5lp88a7vgQgJ5I4o93jfLRAk/gEkxRtyS8wXeg6OIwUKF
exU6wTKK6l29Fpvf5ujMnvlkHx8u5HAvVde/zPNl/hy3FkVg+YiMIJ+zsQYzy5/AurXRBDZwPvYm
jQGmajFV5cqeTO7CBl6lYR4XxXBMJsHNsk4Cl6oQXLSMjQYAONWKp3LprujE+MerJnk8APkO8Nh6
hu9PMph36V0BZgX+BsbMKikrVu811xS2PA3IfYdqI69UqCAK4M1t3p9IDeEvOIPRz9pO6AGxDy4F
uGY9qU2bRVPonxeKDQLMS1Z/V40fsEFCiF8rHWn3IsC4vGvKS6JczPrAwX6f7zts0X9vFfoSyeBs
oXATku0JEF5oB/usqlpv14arQIgFuKaJjMy1hqrGhDKzYdcvxvSXqKx2ABjHGBWkjIyUJ0kY2uJg
msoX99pkfMnwZEW9+0sq+SG18dMpI9MnCOlNHdI7bNeRdT4kNi3H5gX8lGDO6LLnCofxj+etsik9
lGb20a2jWdU0zUGYoLlaadY40epJzzyqGXN1TyMQvgcZhZrUkvFPCU8RS+7gfg2HyLLEeoy1y1Vv
yusN/mhVRXZMejzf5y4avs3XV/x3uSgHjl0tgGghtKK0loJZaJcVM07JQtF/RVv70/zrS3RLLX+v
2+CcV5/jMXrpsIt9NoTMrDkuIkB8BybRzJ0LizOE3F2BZmy79C74UbyKaQLgSwqPuUCab2uGDkdY
CeGY6+CQ9EPRnl7CFkdX32MgH0ctDWYEHZc2V77UGr0gYBlpbVU6vKa70H2wgF6E1ULe//wocRBu
0yw+RuWk7Jl6He+i3o8a2q0uVCvnJbPvI4l6z5ryVHi1//Tz5CW5nJES1QXExXEVFabWgu6PmXWM
nsWut2O/EqkgqGgASpLpFaC8uaYINMSL1tfnzj3u862N+CyObSvW1KFSB9Zqr4Jn2ND89XUEvNPn
9OB3kWjut9Og0t2OETQurQSpXHBfBLWk9CPwPMmPpTaAw4TQWrtw42V4kfKFrmN9AseyhFiWXQwP
R/lDIY4Gayloso/STSIpcJwx+8TxPR17JE6LwQLH+kRsjP4dtZ6/z0AODwYRQDBCL4uSRcZ2A77i
WJXS8qAf84v6abMB5WJvw1QTJS9zmE5JUENGumfcwb93VRG1hEnPsinJszBxDO8MlWb4lqPisQwQ
Mu+l80nvgA0CUw9PasZSJHmWhoEo5dTnySA3Don3HvT47G4TDmk4OnTByMp2fc2IVf8Xgm/Ip84I
cGjdIIfnSWT00aHh9YnJS9JAIcXXtKT9fBiLp8Dm7TXk8x5/igGkYfWPcl0poszL690P7lwD/tNM
cssmqIbs9R4VTveRdgxjjtnpNCr7WuaskIV57wlrHnE624M5NLjalkfjs9Lx4o0J840j2zp8lAN8
OSTR/06gkB2xNEvOB3wkMrudBl0+jS/KxQh5MleqAcgkPNL3FIpgj/dzFH+RxHIrcjw4czvRJeKr
TsgwFfFzzfUhP2W60SO/MrnLp82EZ0fLXqY8v4ZFjXQ64kEJj+NAxrxGZ3V3z0WAKLh9a+dWQz7U
xBc7d6xfwebNlUQLnJPG0lv0FpQg4od+L8eh3cjqDf8diEAkSeFarh5L4SSNvt5nzyX26xfkfnGV
SG3vhKaDe9UK4SLRwitsIU5qhVXVZDnX1HE1t8++kNNBjy36b2wvV4hYXJ2iv7itAKLN+Iz1TRrl
VzeU0YPJBgY1W71zQ3oxYJMpJraTXuBxEbS7bRXRea0Ri4MuKxJ65qdcIoZ08PF+NCQ3B9MvXXeb
FdBiPKZA3fExAhj/US7ghhEyUbYB62jbNTsRtU+YYv11+6I5kXJbTmf2j/0bg7ELUvP2CIfOwQnR
bBwbnxb6fhjOUQFcIJLmGP2ns1Wh2+U4cIv67CzfSpt21hfBm2rKtSR0UIhSnd4py1jeEN6fCVfu
UiygTIQMFtZxvKBMC9G5gQowIHd62XjYpdvsdXaFOhegk/yGG53k060Sv+qriZYE72QvrPqNbkpg
RuIZChGGvp4trM3y6K+PYOYo199P59+N9BjSOgrfdNtdIy937IS3ezgPs7pbxFtJIqQzGQ72Agk1
umpfh6eCAm42pKWJ4F4bSf8eiBB7tjC2AJH2RdThqYwGz0rVvf11zXkPuln4dj77milZlEU6xjXd
nh7ehrRib+GTSc2hYKpyvjXp2B48KSjujMdm9ZBMiCwbOnLVzG8Ma+7ifkp3qfhg/8Y6zDqW1G6j
JUTSyIy4hRM8iAFYbvKm5Z7wuTxs6RQWeWBHMJBzoq4tVl5/ZW/D/8LDEGZNjAeqaxrW7a2IuU1x
0QXZ/unLt/1XpUtPpaauJ/BtekBmRyQdtdZjWYOSYO7rInKuez62Zf+MzOVztR5kyIYoRyF2kdSF
OM2ec0KdE/uLBFEWU7H/SMYKUYcMocd4LbTUGh7oVJ+L15bMardxDsKForSPQ2OkqOCeuCW4aLrm
GUa58lxl3D4pGIgHRI0N02nAAyCjOmrqWRA7coH1jeN1al33sbxelboLRp+yTeBgA5s1yKxILeXS
GqigvOBfl1UZMQjFJO2jINr8FgRnbr9lMGjgGsXsC9PCxS93q9P5hUimICzetEK4ANL4oqxALS+t
hbIEuCBYiTdZ2pPYlP9BcmhuZ34joIo7aaC6tczcCbzr3/Gc7WPrmgp7KWwsDn7SSVziEkg1Mi7K
g3nAvXcfbuGLaIrpNNyXCOLqan+Rbt+Uio8PRBUm9HUAtLzKRG1kGBIbWkLiX3khbuJc3gkRNcmV
OUo5yVjoX4wuoBPQH/9vGPbVzjBgsBp8V0JOBln03+2SWi+8VxgoOBwLijRISuow7GEJbCT+geds
Kp3AyO1E3QJNe2AxiBj9OVwzDBFKA8BaQNO8ZiDdPTz5jXtyTn88XQI141id7+CVz6Twlh/GHdBC
wPusieYI7B5p2Mc6asxzBSnFxjhcvDaTu1oBNHqIlR60VGwjMut1Fb6dp1Cl2Lgtf5rn8rhyyaSU
3+vmFwl4SgvT/MMJsrnHKU7f2ADhzV9JM6rXi9AmdmmJYggC5lH8Uf4AUduebNdZc9cpbjw4lMmK
JPzD6eauwy/AKV4g4iIhvPleEKkGL0W+HcLrhk9/LQA0Xqt3z6LL8Xx9Z4iuKCM9mWYj5F0BWlfR
oXku/ADGVqXnVfyxTnopOgLAg+ueSnWGI1/+IQjWnatCveQdo7dQh31JOfFdDCpwEhth/hrF/v6W
Xx556OBD7oXEwLS9khdJtedgpkF23rxT8tMLzrSEAApIXUC62r19OsOT+q2nMvT2O2KBI2ZNnL1x
qFs92YKtQybhtEHLh6KzAa8I87wKKgS3G16RM3k4qRjp3PT3xTRveUxDoOEO9fkpYdP6QUswGgDi
wYc5fRMvUL9K7/SEpXhMyeRJRgJLWMGMKdb4WJ8t3JM2IiDc002ewcr6n4FjlqQpW+RP8utOcCzV
qx4+HTfILiTN/hrbzdEkxbpDy+Pk00fGjc46UbI+HKmNbjaYldPORjhNuFVdrq0rOiT6oN5N104p
B/kSfxo8pe8NVh6FHRjQIZYPo+ZlCMaOLFmTzinHcTbjnwfxGxl+y6+4wAlXZxDpsjk78jhhESJS
wGrnvnkzJtTbUVaPtCGs39iwVAA45P/84mTNVKhzmJ3zZaJSGCFwoR0VryX90vutxsxqDC49J7RJ
IKVobsA8JjR4myXgnPbr+3mX84p5kBcfxh5rdjga1wHTxKzRA47SPaS6mdCQNlYCVe6iL1G5YaNp
hsZ5t40mbM0h3vI3gSvFjUwhzOCKaeBEAD5lpzMt5NFv/uzPUoVsdjlHhgId9Rn4SIgQodbLnRXy
i0i84wr7RSJ8fb7KJfqKYu3gnHOi1VeFS6q0aAHfBKBVJGK0K1vq+296gR85Nmjyb5y8l7ONP7Ah
cos+xHjJUf8xGTagfmgW1DrmYK6GXjCKdAJpbslUFkpn8ov7nZ62J6wsAjw4epSwMkFMQlplz4aY
VtgAUI5WHQXnOL9qH4PCJzbFv9BuUamF7vQixMvbgyPF3QXMF3vgMN9xE15ycbRh5AGPY2IQi/RM
M94tg1Y6SP9sIHFonk25ze0lw7TXWCqsC852Hcgty2ANVZjmdMhHDniGkcqCOwJMnjd3UKrMzvJE
W94Erth+UgY6EH7HyTcOFZ0v1P5Za1HIq5LvCaCuHhhfUrc/n7rMiQk/pytlVS3WIXl2KHn0v/Bt
ik5lBZr79icj5YEmTzw2qwVK+XPkGUz4k71aeMM1/liBvWOUdrAvlR1Yzc/UHAzeQJ/StnJ7LpBX
eiQOZF/Otbkz7ZZ2Bc0R+oo7yohKImQl95prPAxOaLI1MVk1h74bWExya1SH7e2huDaPLVc+tRvy
ZIisD01WT8Kl7/guaEp6wMAdUcBbzFY6RFmR5dRqpbwGlJo/wmGWDnjvH9IVlM87Zo8/Nr14Slay
/+oR/4i/dJVEapkWr9+ZukXBfXrbwvt87dbsRvaA3iaah+5D5D7sck46h3n+2XEeJJY4UuxvG3d0
/7dMSLB4gdtWwRepMYMlrGtDjRLv5SiZhpT0xK2wr8ZnT+NhUe7oYYO5uix7gZ3fU6kBMyL6HpFp
kvL7JGZmiMoCEaLQZwAeohdwCNIWpZ9Cgpygs9w/7q0MmEHFz5eIoHXg9lvWkEHzvr0f0xoeRqx3
OQ4JlnIpC/o8x+sn+a/9MBb9/2wvzzBa5rOzGMAB71k6RI2XQIhcX9pLk/yyiettGFE22DyxPLnz
QHrsnPHBNsNfWovssykJFiTRXTwIuo3LzezH7kbY3M84ppc9WoIka0eJIn512k6DolBTusRnXJAx
GNb727pdOtnkuCZbrzOD6tVTWDQtrvkUdO8xVoBh7iNi3gGybq6UcyaPx5NlDBTlDO4YMLuvZQ7Y
IKb95Bz8dHPdFJoGSUYoNFKxPeUoe29NR0wOns61ZdyOadFx4zBHzRg99aQ8/kd5pELI2YwyG9nb
vN8dNp+hI73gCv5zwtd7JiCpsy0q9g6VCytAwU3TiXLF/Xj6ibxb7Jr9rsNMH788lwNZPOtBkdWl
q8naX/4WNHtT8NESHtfrkUVgXS5Yzw0PT3GbI6K9hNJXhVWytDDmoPaSEIefgqjGk7tbKWCNUHtm
MhsnGVEycExzKk1NcCVYYqzYYgzUM2HwYrT/5PF5U6lwd/xZv+6AZMe0U1j3+dEVdS9yY3024TGn
8IwG8lqLJxBNL2rQrvgmsnTJGKB/PV9Ye4dWrrwiBYQNL3g94Fi2C2N6iP4ylDxCL5e/25kNUrEQ
r0wUwBKegn/nveZdGfV450kG5bRrQBSObii1htycGxr1iEaPYWBR2UCR6061wP9JFaphzSysu5q1
9UN0PpfW+ei7DSOZDoGiPtVpoC98ni/2nf8sM5KsRpfrI59M6sRPNMRzdAn9ihykVXUFRq2mzGUL
JQfZgZm1Kwdq6MRN2XyOMotks1ogzaogUrRu0Mz/zE5BBaVDCdKirEJVPGtpRevuqdHwf5X97B6q
1gyKTYjBNscVUTK3mzpTqrYWbZE8V8e4crkTrC9uc3OOkdUZ8/unfiYh1Nm8+r9uqTiuBajkEfr4
IiUVu/jSEeKrAQBtjVPX3TTVDz+MukzyxYT/d7ZCoYq+QjWu+PaFCExnJODLrMmic+MUD252uEzq
SEdGfg9/fwSFLBGMIoqZnxcwHFpuou9TTzDDts2lzzOpjUqtyUMvZSOuek6ku7QZDrt3+SyLZOW+
sw155xi+0p0+u6bxQK7nZwIacQuSz+V3qgYtSPcqfsgueXIYtJhYUXTKsmoxuK9znIQnRUHe6YYz
v0NywgiZaAN2k/9sjWVCdhuT1M46/DYJ2KXW5Qxadebu05saykwt1ikkf9cZrkmXI5CgdmYm3hMp
dM9p7FTdYEJE4m5KBDsHbqnh4zuW7UiyJ0BjCNiNkDnbtCnNtniZQ9TbCZa/2BW52AUwZizfJyCg
ChbE2gwXL6RrAAlxJyVr9URyPLw6R23bvosmfOlUvJjnPoA4FLT14T7tKlJHBPARu34yuyyYnQ+T
tls+F9gCAVhm1ql0wNdXdr/hAqvzu72vv03w7YuKNveZF/l770Uivsjr75C7VsS/RWNv8oNNZWkm
bzuZiGZtAld5c6R+dKcb6Vbr4EDm0sKdYqecXYGoy3GqFInHivmQ/36fT/LWfn3PHFXg5rLN3FnC
IwEYRDHnKUHL3h09JVfvw2M4JXHwvsz4pTEpM09rtI0p8JWRR92MbNMdw/k/GXPOxlbJhdTVSfy3
GK8gambU/b2mO9zSOEG5rC89va5jDgXX+GboGzq+bnIfVDRLikHE6zMdhHXFoatvtr+F0/0qYeML
/Ixy/XmCWkhZRx3wPXmLRAkkFJJiGyJgdWEuJQ0XQaTZKaQ7OAiTqJeZiyFZfJ3W0h3+8UD59PZN
gSgFljLu9wgwMHxUn1h6y/T3yJFa64G+tXjCW9VsAYeTZR7FdS0FE8doeF5VjRyhrj9HAaybMrju
RVpDP79W5PcTbcZPvN5O+IfwfGlDXHA6RZLXEZYbmiLMSnvCft0/SysqsgZecXIbF+S98QBjsxMo
ukIRNHtzdQcFVtFQ6RolSuhZrxTPM1FNqTVM3NR7F+Gd7h0QHCWzehmgg2BLa9UXOZyeVPBsOLa7
lrzDFe+F09kRO0ontxHrrMzmhidT0BF1yZAqIFeRNCOHlF3Fkt/tX+brL1NJsMTOawcaDDbhA5IK
/bbWOlIaWPYTye3/jCsE1cYWvKUYr8unaYNhvipr4bi554GyV9m6O6YXHaQmQosH3DRJTAa+p6Ol
if39RXMM8zYTvE3A+FOT13OpyfVf1JClJe+6fZ1WdWiRyKKR4oC9viLIinHn2HDdLeVzpgkO0SjC
Qpa6oYHWZBlj2bIdJyOnP0tlS8fLk268hMBC2cfiMDUcMraU5MfwXBXCOpAGg1emRT4Ty094gD7K
V7EOtlJ36fnWNNRTHoczllxNfptRxlZPmGFnVxge/YVeD4sMvkJGXs+eGTNdIs/BHZljmeB735KX
29Kj6jDHUKf53eX6Sk0/lhfOmiZW8xIDsJ9+ZgrS5imU8lF6xix+ermSUJsyOwDpyyFl+Vf3jM5P
Q6cC36nGVq/O+uOr1IGaiCyodDXLHoq/CxElpRWNaUSHL2CyRaNAQiTC2RYGgZ5F2b7mGSMII1X0
CQnueS0DlFZ0GcVCCaAJReamFvLzkdCtFP5KQISF1aDyVXUOThwTAkymXryv26VSfwVdjgcvrEEi
V4Xo1UYtzvo7+/ldrQnG5B3Zboy1OwThnTYS9BGyXzsBuYv1VqlnzKxSVIIB+A2DknOZGwZr/fo7
UUE+5+Z2MSNg//7LAnnguC5uPIjW5CHTdgobrfHO1vcCK2JGkrHF1FOTrht2QUaTi7ERuLnrrzYn
UOZRxbP8AiD67UVV0E2CQM8yT/WT/wIdLJHKOueZxuQVQj8ztvFdhNcmy4FoogY9KXpTuh/ymH5P
WInrP2I9z3KCsaYt575NJOsDhqA29Ctq6ybPdghdidVpYKUmPEQYBfoseQsDrl9qhQdlYXM2U5IR
I9nU4WU9fcORhWYxWL/oHMLu1wrBpGQvWYg8ej5hWyFeXMkIRBEb+k0PnRaQk/nFpWxfP2CVSj6z
USOfSIMBlkrR+4D4xg5kAlx9NK8Ds2O5nMxLoxmnFLQCXWPved7S00RVNVzelFS+K4FXQyvkmOJf
22mWVvsey5UiXTpPIz0O+pG9Qm+cZWR4BZozl77sLr+f/1oWd636LNFme8hJz6L8X97JC1N7TpOT
QStYbYTDrNRwUlwhoGxM3k8FAjyVu/nahrcIDrkvi2oql8PeenlZn/bDCJjlYvLKHfWP7P6oKEUJ
tdM69ARG0n1Pxy480mYiJ/QwXwOvwRkBOgcJIg82puRBp/RSENR0On9oqySxFKzKd4+9u6rfeyL7
T2hK13a5aLEwbPspZJ0sGsKhx+MFDGPdin/aodOydLFb296vql8TRjz9kdeGQw7I2B/a9QzkdYpY
9VxcOBQ7rGYkGO7+Ka1hg7yEjsOrAPFjYZgwaByBzHOurCIoGNPkjNf07cuCqGG5zks4C5xtOWPY
XT3Ys8SAd9bsIWZaDoZehFdKJpTIWIQdF5FgDKtMyZvZky+WgfMpR4oHnoB/Uax+GDFyjWK1ufPZ
1JMjPpdBgTYYb3v/8nZXm1fksw0nGi/LjUF8kUElMqoyBLcBZn8RVgIMo90jGMrWc5g/Ssf7Q09C
koXqcJwfNIB6hU8TokFN20xYt/yEMiG6A7KzUDima/39SlATu+OQlrDE3f/6I42ZKVAN4EMd70Vs
RyS5YGVVq7tNJl3hewG1nkZUTe13uowXEoxB4X/6bmuBCPrtbNT9taYjBlBdE8OFDJuKLX1iXIdE
3CGHpKrJNf2I5Jd8G8VeRpqMuB5qO1wb9oNNqGMrwd2udGLR3BW+2YndpCD5ECPv3d7oi1xfDjMI
ZvWJj+T/HTrsYXRehLOpTGUIXaW0u21CF+/4XzhnxYZ9A/N/d9DBslo2MZbXHISFTGzYHgqqqZ+n
y9OSb/i/ZNmJNgWsN1nHPLnC8VroCR5gWwsm8HD9E/PZtyfWWAKXg+zzTVoqR3x76/vZMPa0WijE
bjyGhqJ4rn8j8srDo8vbN1kqOiii7WpdQn9C0e55YEGfNCvvflsVUIH7Fi8FOxfdrTYat3Tx9mko
0zPWs74atVkzk0ihDjhEPoKej+PMHhFkEap2U/Ew3dEwh+nKWifcTNBVlogeDTQy5UO1trXE06Ct
f7+jyOHdilRZQ6x+4AHDtt4/fnDQTiQXr+WAeDBrNLU9MJmK4xmMdU+34hi+ZeeHGgpFeiOEoPMp
b2u6BOVjkXERokavUWfDjF+ZsyL6k9NInqTtLO9eVYv9Uzq12iw5qWz4ViCBTfpgPp+owXy3P3vI
QmUGO2+XBI1GLAqT58esUa7Uqe6WYLXVJ3qhUMCBEZrUID+N+uD6PVMYyR2/7uikiFXptulRDx13
UEa1+1WmOAPDxAcLa3xsJKVnHSvwEymObywFFUr0C+It/QTSNSe2aU/Y/8wUO5f89u03SNdbJJ9g
0RZcpR04cL09j9UnFyqui5XLtoeP5wrLeEFrZ3NEqizbdgBC9q+lzXnLbVWmKrOX1AnC/SYGPLmN
ICGA/izmT00gNACDHI2wPNr8FfHUDNnFCvL5bEryhYpPOXVdNT7ytvjhF7/sTAcmRz/uWi4pqgmW
Lpry8O5rtATOH862mYUL89GnMtyQKh+kcYt0Nh2P8a5+zfhZs8ObIcuGE4bJUmo1LfLKJvfTbFvF
cMpkVV+1jJ9myRe2VzrPlzQYU6ZjLVfYec/qI0+4daqcXsl9Rr1GSqEhn2R1PQ+e41nTMU0uirst
Q0J8xW/l5EqteoRi8paLSw+yXND/ZJsJfxnuZedetsEsKaNRleysI+NpBdylPjw9IMB2xmUUySjS
dfSVGvCn3TcO6eF0N7RvUpBxSo5FreiRjChesBg27eAjitCA/DNtxjTiQtq71FYHgyQUS1yPOcyS
1eEUVuJr2tUzBNtjW8N8NHLkVWE43+OdFT/1atO//+baqWB8t15acBeqdf0ySfaAeFXAir/JMBOj
qEvC1QSZW1CF+bYxNo9Z5CRC0H6NTKDEdn7vOMCvagMTIKL4htMb3m/6Y7gT5wiWEPBwQMmfaFfX
eGHa86A26aBJbUbe+9Dys0ZPbFErV/VWD5L5nGkQMCzRIgsRh2t3PbK19pL3mJpCXaNHrqT8wyfK
Ed4KLrVdgjUKerC9pyRZqruq+dSMMiqC95OKKHzw9S6bJJQ7GH9GbDIqURDmLQ6TaoqDNCvUs72/
YzBbEnWcfMuHXbifHC57zEkmzr97/aMOO/NSXIcb/pI26KSokEfZDEPBxEYJUkhIi/Lrpi3EXjhY
1Eso8DBv0W3JNRtow/tOQJ6JOxMweHlBVeZNxyvRB0QMx84CatUlFyptNtDXstTD9UNFNzcMme6w
lkpUggDMFMhhg6oCAJENSFIRf8k9/2Tk3eqHHHf8Ar3GXqsDg5ukc58I2Q2JN0gEAVUGDL7TSKv/
vHEOxS5oJbTZQeEvNhlw67JRiz3t+v9jDGUsc4MFZTzUdYx2vexovUyEG9bq26kGo8o7iuEpxc2q
/BNdSu0DDsf31QME4aEbAv9cDqTqY61qs30XQoosrdvJ1KcaV0Z4qv58VUu8ip5QSRH3HkDD5m2q
NQH7UUXBWjsWlbOoxukpCNWRqtSnoF4ZAE42EvqNwg4D/RIOf06BMjhOKaOvblRK8NkdWqM/LNNc
5UPcJk/Hu6e0s7FvMfCF/EZUJkLP+cCVh0diwZxUtxVo2kVAVE/ImfxOzZXtJ2//jwsgA32GOsc4
fHgWgCJYNw3IbIWZ0ugPyHlI+zxDushgG9ClmNaGRDs2+ePFFyPiH7W2YMeKhjRmncYNOoIw81jX
uCqftlH45+994OI++Ttwd+GpqFxP8w0U0vwKrULoLnRkwoMJBkDzGTaEdiJr+yz1Af1Hmdn5sopI
W9SBz4xwwsB4QKkKzLdGhClbklAtUjU/zXOoHi/w1kWOvOO/BZuNssLrkovkUIbjpWewch4rDtSL
ac0N0mOeidmbbZz6qvI7MHhaiEONpenSLFAIjvRxwV4jqpNyyZ4eUUURi/5CZSaelBru2+FIlnsO
ScP25upGG18/NrJ8XNx4/zSL8SoLiY/D9tlydytu4KUrJmBlHVb9HWwKXv24Txxls0bOFd6njDyx
YsHqSPmUXRWzd7DM8m4Zj0QTM0bkm72si7F2vmmG2oWLArH1F9XGvWWDTwVZrM7h4EqmBx/PPGCb
9vxHhgYi/Bl2l+xBQAe4FnWNX52hc/VnM1TVC0UEWhF7WE86mXlopN/HUmu56mcAPbk06DxjqE1N
0QMTqyoGiFvL0JBip9oX3hRW6m3fWlL93qmwji3D7hNkuXrm70m0pPiyV2jiQoYjkK8QMq5Oudx6
X0z+LQ57Z6UHCiYp5+73/bVZWpJnx9ukU173y3cV8LbUqzE/Kh4XA1UFNHeQPywgQ7OdDjT+Wa5S
SfD3nJQmtqhbY3M63Zm7zMQhpvp0DDOIDdypmIdfQIUwMcygnwKbCYsZbXRtPVne/gJ6otm5iDAv
bt25WjcJAIVyu6aQ3C8Mut85O0MABvU2eTHKmMDG5K6U1uDKRYmQ3QlKuEcFzUJDJ0STm3sWAdfn
aij4XFsos4YGTmzlWRTDvTGm78iZsAaPHuq45H8+Lp55g6zRd+IJ3twHwksXXveW005ZPx6rNdoU
nw52SQs2Amor7PwjKhrqcIWtIktZzQaY1UgRkYk3G6gO63D3kPaMq8JKt7tH2LtTt8Y9IhsO7xFM
DBLREQtjqilGQliS1N9WXPwjSCf3+H0afq4lEmX7ml6fWic8Ow8XpwsNUnDkE5aK/KKpi2UEsrq0
yG8A4FnsIPawAan1icELyNSHXtBDFKSL+Vwpv5Bwuk9g3x0uxSJ/+OntI3L/ts8BAr3E3dtOgWp9
B4vxImIWNZdgtmTOZ1Ro7AWM6hAf/jTrwX8IEPBMrUyX3h0p9wZCn3iNWhRm1G/q+FmlqiiTtkvJ
lzktB0tLg/rJHBqTkK0frRefsRp9wt6ZxIsVB0rZxgK4MfgmMNpFc15Hxhf7oZF/uhnOu+zmfFvi
j2Zamw44RASX0Fb+iyC9uJU+jl9JLx18JD3oFGQeU1h2796/VSzGMdufvVdgKp0aXfrionGBpUyE
bX3uM0SyutuDcgnNV9mHy6BLc9MxwSxcBTmZIKEESk9w6BFi+OT0DUb5PyntrQsXIvlZzLN4+Ogt
xkdpvrD/NhbSs1zn6xMRPgNlLyZAxVttVQ+qLW1b+IaRKnr4UiDM6JkXlF0yHRWkS7YKShVhEeSD
wApC6ND/eqwtVt4HNU659FGb7sYBSalt80cIsm9CZDfUNIFYkFh12COBZPlD/EuHc6K2Q8lO9Lqc
xm8o4zhAllZGzSZRV4tnqnbVOJeFjhcgLyOXR3dtokT94CjAOThNkAnPgUxiDAxkNccEDMShllXf
UnbDE5XTxoZzYj5TJUuC5wPrZNuCk1Iw9p1Cfz7pJ9tzGL3rrldUvxqeVge9TDjUE3pZk1SEhsXi
1F2yUKpwRSp12RmSPb30y9NQ9UGMphuuEVmmufy70hNYXEXF8wIX8b4LMt2ngCM9e4BTnryrYKz/
8sNp7f/J4Dmcq9w/JC160qIlqcQhY4Xw7L4sJkofePbj001ml27VdmN8OU5/dEc/96wZ1X2DcZZn
G/Ou9gHgtZeFAs70isIeo0g08EV5Ajv6ScOIrjQZ1H+7sULhSmd2wN9fjI5awWY9mO3xs+bgXp1A
DQ0m4Q7gtjRytfm+XDiaBq7nVR5Ceez9vOewBEHOovJqijgbm7GWquuv8Oe7A8a1SADr3PB4vEa0
/ZBHccbDKaWQv1bOYNEcmGtd+4c1bIT4k66Tj2Ugh1vGODLSVob76PvFCgCQzIKp9Wks7hbPHAL3
vCjblDJxTgNE2Jv3n/4wadE8nItw3BVeF5fJG07sLwsI8CzzCfb5qTmg7Qpe0S7RkSdqLzSVTKBN
+LXI2M1FiFBY1VbbuZFMhasg9n9wv+k8hRg42jKY8TjWhj+TdXrY9OTLwgRK+qYU/o1om81/NmdG
XwlIUq7AvwcabLySo7jp1eEgvdnZ7Y4Lz5+ld5WDcK4Ao0Gu0+Q709aFUnM+wF08xR6JcNNiPIBc
V/FMP5lX6ysYD9vvyyqqKOa/0Lr8wSr3kdfTM8lBufL31cBtJlypPUmbS/GYFbOSCDZzVMQswEnB
WgREhfTPwzwKxZNJeVwsdh6EbE13/pXGggS1IPXNBSenm1xYGkUABeH3TA68KQXslt+GtU4/mDjZ
Ql+ZEIkGzIOHS0CIwd79xu28oieYMK2LvM9sCvR1R/ox7xcmsBGdlThJgTkAJTb7ApBgCCD2gqMf
j8X8jL5Sw4vpy5BPUfI1SDxOhCUSzo+mX8Kb/B/m0mjL7xMRihY3h8Otv6+QI4bykJcr6UXQEE43
iC9sNzvgVonuEKEY6uL4BGPI6ol0Mft2m0+mCDQMKSA7GCUYQ6+YYgoeqSehGim5IMwAjPSwwXxj
Cwtk+Uecu1l4j3yI/GG3K86G/SlYUsdL8/cuKXc8xodFcmHcGBKUZqxA/7UA0UWZG9bUbC5dCLHg
jgfrRkLjQe1aTw0HiUniIC/Aoe72Jblm/ki4PgGYZPaRIT/Kz5LmJy4TV/37mjDtCKXam3Uyk+0u
us43u1c/rVYWZk0IotSUCM14N0ynFla/AueT6qKzBdCTUdU79yH3oA++F245mxVu5ojVHwtrSmEA
yadfZ2AkYRuU2jiam29GxUobgimMUwuAmjZIw6lNVuAXnLMV7TBu2bcb62HBwM8J1UOouOf6S+Qe
Tb+W2/6csa1YfPDo3BZmL38dADvHJaqEpFYl2AtXQymmd22RNi7CQSJHyGOlhYLnd+9X9NrBJohu
BsdzSe9P7V+9Uj0ak7t4ZvPONPE0IDCQj+mBqMkkX2fC2EWRpnYc04cMFvAIO+punhCsHQA15Zwt
VzD7nZHR9aww1ITElxYfAnB9f5/k26WI/pBXatllt/Ev3tAa3EaL8YJoOZIR7xC/fzz2oydg7yBR
Lig9WDyj6GQ2Bv6n2kquYskLhtEtPjkvh6VCWuoH8VTDx95mH5QbfUw1B12s6T0n7KT2n4TEYo3Z
WkFD3MiZVJ4PNQ+GbpedKovhfRYoFU6VobXCb5edaA1c2w6QwRLs11RuwRIwleSFK+AgZ1frBjGB
mxr1soMsMSMoY16R61oLf4ojSIZMkXQsSwm+6h1nD+3TklPD4ELRxLHUavOw8vvvhyRG34GGIP34
cJ4Agm/5KUO7PJUCzyJ12qbWXhSzlsIqxK+/OjHzH/78DLWfAEnMkTau/WJxm58WqeK+mnFSU65Q
ytwxUz9xWyL4tugCs2MxjYr5ahUFsnjS0B5ZRVf65PHBEGKt2upiO7brI1XD8B5Kz1QmaxlBU5rK
PX0YpoUdcr0YuBN1WXrtEZRb9S55ocHPThkPuID055OXJtw9g3z74ywEb/Sh5Fxi5jR11xC0WAdq
zni89YWL8OeIwONY7eMHamrEE4lpkxz2Xq2tSqiCQLNSpbocQOQjiSdRhi6Zba5tSAS7MPoLPa+P
RvvZAzCAlzX5qPZVkHZUtGUzMOXkqAlDLHguCnBPipnud75pN2Wcw8BeEP6QHVQV0OBYVfg9DRLU
+UjCk4v0Qr57sqH90kPBJg/OuLe1l7mDQ6UbT333+4Xkklh50noKSWi52xPvvm6OctbgEWjilk/O
XYebinl/5nm3R7wJE9YxO0xsP4k88A6xYxC1FdrEh4g5QpgIRGm9kd0SqZziWDpdkLUTA1pW97W0
yzUxNllCKHjv48DaoEkNMg58HoANASm8ZueVgnMjpomyL81EOZfT1DXkLlmxuQrJk2YUxs5hft3w
fFyBOHb5uL61XIN6ZsBJ+50lIkbIUGsod+L2BySyQNbWILMg38eqbbbC4TrIXg2myYPXB+43uSbp
fIERoycxiMXaJTJkC2wl6ZkhEH5ujuXUXyOM9/2oHNgcdj14SC6Po4OKld3chJICbAQT2VPsq8wc
y1PJxg8JO+MKZg3mQ2lmyJhIPf6LwoAXEoU6/yW7dXdbH6HL7SflZJJaE16dpOvTNCv7nplc9V3q
30kQuqmnIhrbrxjwEjYau610EsOouljQFTaAg0scqWSuWKdGNcDdv/HZgg9hhtBk6FNUSNhtsCQU
TpuLjJjzl8+b6Z+KrZhEabBRRGLoFfDwGmFpJbCv2PXKfyi7IJd1rxYzl4bbOFThYgv74q38a0K/
JlNO5tO/EWhEEwHun4iCv4tLWtZeE/O5WYwKMbIgUJX2315zFNBWRhBFVxMMCPKp9oQoXSZCWTeI
CkAFZhfQFm1cEzZiGtMZa6A32+CsFABtcFjdg3P1gUtHIHBWvTNkXcvJG7BpYppCbYxMPwdOIYuo
lwb7i2QXwbvONZXxkPoQKmPCKYs5WnVmyCh12TeaP0RGHvE6Zs9JCzvbwGTimibeT7xjf71vXtnh
Wub5Nj3QRnJoXiXPls6Pz5YmvRLofqJoLVSKZ5QE/dvtWRX4solR2W/WbTqpS8D3GmdomPqi5iy8
PEgV+/6GA4YKXl/ll+3pW/6p8kw0lyc2Mgg2HtPHQDrypE3WINlIEAaJn9ZojTNdxsxgFrCPBu/1
bULhLNiCdPMa+An0ohs/8yjKgWZjENzDUHHdFOM26OXuIZ6IS1f9+Fz41cfJTp5Nj/PKxHNSGiY5
cp9WDTJmGpNtiS5TWDIUjvUONevCWK45PsyVxmOfmh+HTp8exCeJAladYfHfcXGP4LY6x6Rv5qC7
8HcylIMGMiLfrab2Dlx1fXabm54JVW1QRNxGZVps8siybmOiqJuDbOVJG7QnTd0cEJnSaC9F4EIl
wFMaBV/+oS3rTdJpp5vWH0j8xy15hvMUPe2XphWUg+ab4O+0FKkRwJzE9pYHgjGSzISjynaES7sG
oqbYLfNO36f3yWO7dcF4h2+aYPp79Gsz+NmgDbyV22fE2gCDkV9tMLAfx4YuDTRAqWJSL+gROI65
JWlDYicVqRB08lByZklDTkWsmvgnU/FU9AfJ7Oaov9prsSbMxzJazvXHyVxb2eyrKqbkuaMd4F5B
bBA2AoWXCSPYekhsJkmKecJQTZp9MyTAmApr9/54IU6J8fH67DGFEjCKLlfxZVnWhsmS9PJ35Isq
RxuQK+AWd4lkHrI1HphBZ7y+xSw3qZLiOg63zWTAFB+ixmcwzt1mubNP1OiWePrJm3vComS2ueN4
2WlIpDzRxgoE2qEPQ3CIRtB3I9e6abuU/CRUg5vpkXnVY/iPCJFX8Y2BNcorT68KC7QtLRKDpNLR
fsTS0d/tRVQIL+SXPAmkM5oi/l3WeBswQgQbH5iXt4M51LX/95q/iaXbWqNkiWDfS4cx5eLOCQq5
JKyIrdwMORGbHHSCd/w0A+xI3KwGluHC6VcuhPjgj247aLdRinAJ8u3SB4V0AARxvZrIdYHkflfU
YB5l/dOcfd37G9enkWLRVq4OI0IVb8LcJSrvDZZJ4fAY7KClQ9+W0gx3OYsdkZWkMgqQ5vDc2/Ey
WEQ8aplX8ALhD5KFNZfyPcnll5Uv8/g0rXmG3UxWFGzf70LQ+HELt/yN00Fvp/mOcpdLjG/6q0Uy
BWptrynAWyBwRM40tdJTAawrM3QNXRbznufGEWXZ8rIAj49ocPiiCfb12rtx2gp+L3Q949QJM5kc
BvsbT0ATUeVKzd1qXqS8L85oUpTOcRAo0eZLNV9GOzb2+hk21koiGUAxvM5KnorSrdTU43Og3625
kBTdUXUHg9+Sbby3BMaBx61/rH1nD9UHsYIIIlfrBMJxzgSce53mWqM4zT81qltUdrPko1jXJc+B
XTWnSAQko+QDXXmiC+SRCDMqPxxHlzHWqpUpOpZRialMGy/u07ZkZKihe00MQXiUR6Ittw8f1D5X
3t8mlpCdmKmOYZC9JaN7fs+8/yrxKffb5N4OAvwPBDsS6xQVmCNP3ZU8U4RXMEr+u+tw7WNsyX5S
y6ap/WoxI3P3vCJJDKFV0eTG6JOopLJv43x44Ue9ygXC7CdU8MsghGC2RXuZOwbhL52dHSpLeFZm
c+kcZxGAoGERuMPY4GQYy98hxWTvB01FuP2UhS6ETaYCo6peY4tRg20L21cT4GDqU9YUYBDyDqsE
MXWB+pj1gZ+UrRe8rDXEJCkJImBhdPAcXDL967sB8TV8uevVw0RByn1MPilnfrW2L5EVvhohqbIT
FoMJsPZbo/ZvHsCHgqGi8TdBlDAshfTlRTzXSfieZ0zEfMivQrPXHfMmi/kd/DcIJmSUvUEjY8Sp
IcmO8qdMBn43J9WPvOgppj40xV7Cr8WIKLHN7MjpqrA5huHWWZb+SZtNXy8U8kPotjfnXllM07+o
LPKDuWoVVyca8StljsS4Q6Z08lqQ3vIBl60E3CNeBkJaJhvV34xkTtpdwufTn3dL9YoAr/aR9uQi
1SZAlRpjLG4lj+Tio91HEKIuxFD3jqD+GvBkhvVuoTehhL2Tk1nmDE1YNykeNTrBKStghn62xtIJ
PzlTd8GaCVrmHf3NMd4nzxYMTdbru6WOvUvRvJQCMEL1BJBQaRID5sEpvFG4sL4yMYcy/YibhoAX
QmFfkzQY
`pragma protect end_protected
