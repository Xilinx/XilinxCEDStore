`ifndef DMA_SOFT_DEFINES_VH
`define DMA_SOFT_DEFINES_VH

`define SOFT_IP
`define KESTREL_BASE

`endif
