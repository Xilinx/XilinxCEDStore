// ////////////////////////////////////////////////////////////////////////
// Copyright (C) 2019, Xilinx Inc - All rights reserved
//
// Licensed under the Apache License, Version 2.0 (the "License"). You may
// not use this file except in compliance with the License. A copy of the
// License is located at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS, WITHOUT
// WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. See the
// License for the specific language governing permissions and limitations
// under the License.
// ////////////////////////////////////////////////////////////////////////
//-----------------------------------------------------------------------------
// 
//      PCIe4 Model - Core Top
//
//-----------------------------------------------------------------------------
`timescale 1ps/1ps

//-----------------------------------------------------------------------------
`define PHYREG(clk, reset, q, d, rstval)  \
   always @(posedge clk) begin \
      if (reset) \
         q  <= #(TCQ)   rstval;  \
      else  \
         q  <= #(TCQ)   d; \
   end

`define AS_PHYREG(clk, reset, q, d, rstval)  \
   always @(posedge clk or posedge reset) begin \
      if (reset) \
         q  <= #(TCQ)   rstval;  \
      else  \
         q  <= #(TCQ)   d; \
   end

`define PHYREG_EN(clk, reset, q, d, rstval, en) \
   always @(posedge clk) begin \
      if (reset) \
         q  <= #(TCQ)   rstval;  \
      else  \
         q  <= #(TCQ)   en ? d : q; \
   end

// Fast2Slow
`define FAST2SLOW_MODEL(bit_width, rst_val, mod_name, fast_input, fast_clk, enable_input, mask_input, slow_reset, fast_reset, slow_clk, slow_output1, slow_output2)   \
   xp4_usp_smsw_gen4_fast2slow #(.WIDTH(bit_width), .ASYNC("FALSE"), .RST_1(rst_val), .TCQ(TCQ)) mod_name (.fast_bits(fast_input),  \
                                                                                              .fast_clk_i(fast_clk),   \
                                                                                              .enable_i(enable_input), \
                                                                                              .mask_bits(mask_input),  \
                                                                                              .mgmt_reset_fast_i(fast_reset),  \
                                                                                              .mgmt_reset_slow_i(slow_reset),  \
                                                                                              .slow_clk_i(slow_clk),   \
                                                                                              .slow_bits_ns(slow_output1),   \
                                                                                              .slow_bits_r(slow_output2));

`define AS_FAST2SLOW_MODEL(bit_width, rst_val, mod_name, fast_input, fast_clk, enable_input, mask_input, slow_reset, fast_reset, slow_clk, slow_output1, slow_output2)   \
   xp4_usp_smsw_gen4_fast2slow #(.WIDTH(bit_width), .ASYNC("TRUE"), .RST_1(rst_val), .TCQ(TCQ)) mod_name (.fast_bits(fast_input),  \
                                                                                             .fast_clk_i(fast_clk),   \
                                                                                             .enable_i(enable_input), \
                                                                                             .mask_bits(mask_input),  \
                                                                                             .mgmt_reset_fast_i(fast_reset),  \
                                                                                             .mgmt_reset_slow_i(slow_reset),  \
                                                                                             .slow_clk_i(slow_clk),   \
                                                                                             .slow_bits_ns(slow_output1),   \
                                                                                             .slow_bits_r(slow_output2));

// FF Chain
`define FF_CHAIN_MODEL(chain_length, chain_width, rst_value, mod_name, clk_i, rst_i, ff_out, ff_in)   \
   xp4_usp_smsw_phy_ff_chain #(.PIPELINE_STAGES(chain_length), .ASYNC("FALSE"), .FF_WIDTH(chain_width), .RST_VAL(rst_value), .TCQ(TCQ))   \
      mod_name (.clock_i(clk_i), \
                .reset_i(rst_i),   \
                .ff_i(ff_in), \
                .ff_o(ff_out));

`define AS_FF_CHAIN_MODEL(chain_length, chain_width, rst_value, mod_name, clk_i, rst_i, ff_out, ff_in)   \
   xp4_usp_smsw_phy_ff_chain #(.PIPELINE_STAGES(chain_length), .ASYNC("TRUE"), .FF_WIDTH(chain_width), .RST_VAL(rst_value), .TCQ(TCQ))   \
      mod_name (.clock_i(clk_i), \
                .reset_i(rst_i),   \
                .ff_i(ff_in), \
                .ff_o(ff_out));


`timescale 1ps/1ps
//-----------------------------------------------------------------------------

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_model_core_top 
#(
     parameter           TCQ = 100
   , parameter           KESTREL_512_HLF = "FALSE"
   , parameter           IMPL_TARGET = "HARD"
   , parameter           AXISTEN_IF_EXT_512_INTFC_RAM_STYLE = "BRAM"
   , parameter           FPGA_FAMILY = "USM"
   , parameter           FPGA_XCVR = "Y"
   , parameter integer   PIPE_PIPELINE_STAGES = 1
   , parameter integer   PHY_REFCLK_FREQ  = 0
   , parameter           CRM_CORE_CLK_FREQ_500="TRUE"
   , parameter [1:0]     CRM_USER_CLK_FREQ=2'b11
   , parameter           CRM_MCAP_CLK_FREQ=1'b0
   , parameter           AXI4_DATA_WIDTH = 512
   , parameter           AXI4_TKEEP_WIDTH = 16
   , parameter [1:0]     AXISTEN_IF_WIDTH = (AXI4_DATA_WIDTH == 64) ? 2'b00 : (AXI4_DATA_WIDTH == 128) ? 2'b01 : 2'b10
   , parameter           AXISTEN_IF_EXT_512= (AXI4_DATA_WIDTH == 512) ? "TRUE" : "FALSE"
   , parameter           AXISTEN_IF_EXT_512_CQ_STRADDLE="FALSE"
   , parameter           AXISTEN_IF_EXT_512_CC_STRADDLE="FALSE"
   , parameter           AXISTEN_IF_EXT_512_RQ_STRADDLE="FALSE"
   , parameter           AXISTEN_IF_EXT_512_RC_STRADDLE="FALSE"
   , parameter           AXISTEN_IF_EXT_512_RC_4TLP_STRADDLE="TRUE"
   , parameter [1:0]     AXISTEN_IF_CQ_ALIGNMENT_MODE=2'b00
   , parameter [1:0]     AXISTEN_IF_CC_ALIGNMENT_MODE=2'b00
   , parameter [1:0]     AXISTEN_IF_RQ_ALIGNMENT_MODE=2'b00
   , parameter [1:0]     AXISTEN_IF_RC_ALIGNMENT_MODE=2'b00
   , parameter           AXISTEN_IF_RC_STRADDLE="FALSE"

   , parameter           AXI4_CQ_TUSER_WIDTH = 183
   , parameter           AXI4_CQ_TREADY_WIDTH = 22
   , parameter           AXI4_CC_TUSER_WIDTH = 81
   , parameter           AXI4_CC_TREADY_WIDTH = 4
   , parameter           AXI4_RQ_TUSER_WIDTH = 137
   , parameter           AXI4_RQ_TREADY_WIDTH = 4
   , parameter           AXI4_RC_TUSER_WIDTH = 161
   , parameter           AXI4_RC_TREADY_WIDTH = 22

   , parameter           AXISTEN_IF_ENABLE_RX_MSG_INTFC="FALSE"
   , parameter [17:0]    AXISTEN_IF_ENABLE_MSG_ROUTE=18'h0
   , parameter           AXISTEN_IF_RX_PARITY_EN="FALSE"
   , parameter           AXISTEN_IF_TX_PARITY_EN="FALSE"
   , parameter           AXISTEN_IF_ENABLE_CLIENT_TAG="FALSE"
   , parameter           AXISTEN_IF_ENABLE_256_TAGS="TRUE"
   , parameter [23:0]    AXISTEN_IF_COMPL_TIMEOUT_REG0=24'hBEBC20
   , parameter [27:0]    AXISTEN_IF_COMPL_TIMEOUT_REG1=28'h2FAF080
   , parameter           AXISTEN_IF_LEGACY_MODE_ENABLE="FALSE"
   , parameter           AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK="TRUE"
   , parameter           AXISTEN_IF_MSIX_TO_RAM_PIPELINE="TRUE"
   , parameter           AXISTEN_IF_MSIX_FROM_RAM_PIPELINE="TRUE"
   , parameter           AXISTEN_IF_MSIX_RX_PARITY_EN="TRUE"
   , parameter           AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE="FALSE"
   , parameter           AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT="FALSE"
   , parameter           AXISTEN_IF_CQ_EN_POISONED_MEM_WR="FALSE"
   , parameter           AXISTEN_IF_RQ_CC_REGISTERED_TREADY="TRUE"
   , parameter [15:0]    PM_ASPML0S_TIMEOUT=16'h1500
   , parameter [31:0]    PM_L1_REENTRY_DELAY= (CRM_CORE_CLK_FREQ_500 == "TRUE") ? 32'hC350 :  32'h61A8
   , parameter [19:0]    PM_ASPML1_ENTRY_DELAY=20'h3E8
   , parameter           PM_ENABLE_SLOT_POWER_CAPTURE="TRUE"
   , parameter [19:0]    PM_PME_SERVICE_TIMEOUT_DELAY=20'h0
   , parameter [15:0]    PM_PME_TURNOFF_ACK_DELAY=16'h100
   , parameter           PL_UPSTREAM_FACING="TRUE"
   , parameter [4:0]     PL_LINK_CAP_MAX_LINK_WIDTH=5'b01000
   , parameter [3:0]     PL_LINK_CAP_MAX_LINK_SPEED=4'b0100
   , parameter           PL_DISABLE_DC_BALANCE="FALSE"
   , parameter           PL_DISABLE_EI_INFER_IN_L0="FALSE"
   , parameter integer   PL_N_FTS=255
   , parameter           PL_DISABLE_UPCONFIG_CAPABLE="FALSE"
   , parameter           PL_DISABLE_RETRAIN_ON_FRAMING_ERROR="FALSE"
   , parameter           PL_DISABLE_RETRAIN_ON_EB_ERROR="FALSE"
   , parameter [15:0]    PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR=16'b0000000000000000
   , parameter [7:0]     PL_REPORT_ALL_PHY_ERRORS=8'b00000000
   , parameter [1:0]     PL_DISABLE_LFSR_UPDATE_ON_SKP=2'b00
   , parameter [31:0]    PL_LANE0_EQ_CONTROL = PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505  
   , parameter [31:0]    PL_LANE1_EQ_CONTROL = PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE2_EQ_CONTROL = PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE3_EQ_CONTROL = PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE4_EQ_CONTROL = PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE5_EQ_CONTROL = PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE6_EQ_CONTROL = PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE7_EQ_CONTROL = PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE8_EQ_CONTROL = PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE9_EQ_CONTROL = PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE10_EQ_CONTROL= PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE11_EQ_CONTROL= PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE12_EQ_CONTROL= PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE13_EQ_CONTROL= PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE14_EQ_CONTROL= PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [31:0]    PL_LANE15_EQ_CONTROL= PL_UPSTREAM_FACING == "TRUE" ? 32'h3F00 : 32'h3505
   , parameter [1:0]     PL_EQ_BYPASS_PHASE23=2'b00
   , parameter [4:0]     PL_EQ_ADAPT_ITER_COUNT=5'h2
   , parameter [1:0]     PL_EQ_ADAPT_REJECT_RETRY_COUNT=2'h1
   , parameter           PL_EQ_SHORT_ADAPT_PHASE="FALSE"
   , parameter [1:0]     PL_EQ_ADAPT_DISABLE_COEFF_CHECK=2'b0
   , parameter [1:0]     PL_EQ_ADAPT_DISABLE_PRESET_CHECK=2'b0
   , parameter [7:0]     PL_EQ_DEFAULT_TX_PRESET=8'h44
   , parameter [5:0]     PL_EQ_DEFAULT_RX_PRESET_HINT=6'h33
   , parameter [1:0]     PL_EQ_RX_ADAPT_EQ_PHASE0=2'b00
   , parameter [1:0]     PL_EQ_RX_ADAPT_EQ_PHASE1=2'b00
   , parameter           PL_EQ_DISABLE_MISMATCH_CHECK ="TRUE"
   , parameter [1:0]     PL_RX_L0S_EXIT_TO_RECOVERY=2'b00
   , parameter           PL_EQ_TX_8G_EQ_TS2_ENABLE="FALSE"
   , parameter           PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4="FALSE"
   , parameter           PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3="FALSE"
   , parameter           PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2="FALSE"
   , parameter           PL_DESKEW_ON_SKIP_IN_GEN12="FALSE"
   , parameter           PL_INFER_EI_DISABLE_REC_RC="FALSE"
   , parameter           PL_INFER_EI_DISABLE_REC_SPD="FALSE"
   , parameter           PL_INFER_EI_DISABLE_LPBK_ACTIVE="FALSE"
   , parameter [3:0]     PL_RX_ADAPT_TIMER_RRL_GEN3=4'h6
   , parameter [1:0]     PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS=2'b00
   , parameter [3:0]     PL_RX_ADAPT_TIMER_RRL_GEN4=4'h0
   , parameter [3:0]     PL_RX_ADAPT_TIMER_CLWS_GEN3=4'h0
   , parameter [1:0]     PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS=2'b00
   , parameter [3:0]     PL_RX_ADAPT_TIMER_CLWS_GEN4=4'h0
   , parameter           PL_DISABLE_LANE_REVERSAL="FALSE"
   , parameter           PL_CFG_STATE_ROBUSTNESS_ENABLE="TRUE"
   , parameter           PL_REDO_EQ_SOURCE_SELECT="TRUE"
   , parameter           PL_DEEMPH_SOURCE_SELECT="FALSE"
   , parameter           PL_EXIT_LOOPBACK_ON_EI_ENTRY="TRUE"
   , parameter           PL_QUIESCE_GUARANTEE_DISABLE="FALSE"
   , parameter           PL_SRIS_ENABLE="FALSE"
   , parameter [6:0]     PL_SRIS_SKPOS_GEN_SPD_VEC=7'h0
   , parameter [6:0]     PL_SRIS_SKPOS_REC_SPD_VEC=7'h0
   , parameter [1:0]     PL_SIM_FAST_LINK_TRAINING=2'h0
   , parameter [15:0]    PL_USER_SPARE=16'h3
   , parameter           LL_ACK_TIMEOUT_EN="FALSE"
   , parameter [8:0]     LL_ACK_TIMEOUT=9'h0
   , parameter integer   LL_ACK_TIMEOUT_FUNC=0
   , parameter           LL_REPLAY_TIMEOUT_EN="FALSE"
   , parameter [8:0]     LL_REPLAY_TIMEOUT=9'h0
   , parameter integer   LL_REPLAY_TIMEOUT_FUNC=0
   , parameter           LL_REPLAY_TO_RAM_PIPELINE="TRUE"
   , parameter           LL_REPLAY_FROM_RAM_PIPELINE="TRUE"
   , parameter           LL_DISABLE_SCHED_TX_NAK="FALSE"
   , parameter           LL_TX_TLP_PARITY_CHK="FALSE"
   , parameter           LL_RX_TLP_PARITY_GEN="FALSE"
   , parameter [15:0]    LL_USER_SPARE=16'h0
   , parameter           IS_SWITCH_PORT="FALSE"
   , parameter           CFG_BYPASS_MODE_ENABLE="FALSE"
   , parameter [1:0]     TL_PF_ENABLE_REG=2'h0
   , parameter [11:0]    TL_CREDITS_CD=12'h1C0
   , parameter [7:0]     TL_CREDITS_CH=8'h20
   , parameter [1:0]     TL_COMPLETION_RAM_SIZE=2'b01
   , parameter [1:0]     TL_COMPLETION_RAM_NUM_TLPS=2'b10
   , parameter [11:0]    TL_CREDITS_NPD=12'h4
   , parameter [7:0]     TL_CREDITS_NPH=8'h20
   , parameter [11:0]    TL_CREDITS_PD=12'he0
   , parameter [7:0]     TL_CREDITS_PH=8'h20
   , parameter           TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE="TRUE"
   , parameter           TL_RX_COMPLETION_TO_RAM_READ_PIPELINE="TRUE"
   , parameter           TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE="TRUE"
   , parameter           TL_POSTED_RAM_SIZE=1'b1
   , parameter           TL_RX_POSTED_TO_RAM_WRITE_PIPELINE="TRUE"
   , parameter           TL_RX_POSTED_TO_RAM_READ_PIPELINE="TRUE"
   , parameter           TL_RX_POSTED_FROM_RAM_READ_PIPELINE="TRUE"
   , parameter           TL_TX_MUX_STRICT_PRIORITY="TRUE"
   , parameter           TL_TX_TLP_STRADDLE_ENABLE="FALSE"
   , parameter           TL_TX_TLP_TERMINATE_PARITY="FALSE"
   , parameter [4:0]     TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT=5'h8
   , parameter [4:0]     TL_FC_UPDATE_MIN_INTERVAL_TIME=5'h2
   , parameter [15:0]    TL_USER_SPARE=16'h0
   , parameter [23:0]    PF0_CLASS_CODE=24'h000000
   , parameter [23:0]    PF1_CLASS_CODE=24'h000000
   , parameter [23:0]    PF2_CLASS_CODE=24'h000000
   , parameter [23:0]    PF3_CLASS_CODE=24'h000000
   , parameter [2:0]     PF0_INTERRUPT_PIN=3'h1
   , parameter [2:0]     PF1_INTERRUPT_PIN=3'h1
   , parameter [2:0]     PF2_INTERRUPT_PIN=3'h1
   , parameter [2:0]     PF3_INTERRUPT_PIN=3'h1
   , parameter [7:0]     PF0_CAPABILITY_POINTER=8'h80
   , parameter [7:0]     PF1_CAPABILITY_POINTER=8'h80
   , parameter [7:0]     PF2_CAPABILITY_POINTER=8'h80
   , parameter [7:0]     PF3_CAPABILITY_POINTER=8'h80
   , parameter [7:0]     VF0_CAPABILITY_POINTER=8'h80
   , parameter           LEGACY_CFG_EXTEND_INTERFACE_ENABLE="FALSE"
   , parameter           EXTENDED_CFG_EXTEND_INTERFACE_ENABLE="FALSE"
   , parameter           TL2CFG_IF_PARITY_CHK="FALSE"
   , parameter           HEADER_TYPE_OVERRIDE="FALSE"
   , parameter [2:0]     PF0_BAR0_CONTROL=3'b100
   , parameter [2:0]     PF1_BAR0_CONTROL=3'b100
   , parameter [2:0]     PF2_BAR0_CONTROL=3'b100
   , parameter [2:0]     PF3_BAR0_CONTROL=3'b100
   , parameter [5:0]     PF0_BAR0_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF1_BAR0_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF2_BAR0_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF3_BAR0_APERTURE_SIZE=6'b000011
   , parameter [2:0]     PF0_BAR1_CONTROL=3'h4
   , parameter [2:0]     PF1_BAR1_CONTROL=3'b0
   , parameter [2:0]     PF2_BAR1_CONTROL=3'b0
   , parameter [2:0]     PF3_BAR1_CONTROL=3'b0
   , parameter [4:0]     PF0_BAR1_APERTURE_SIZE=5'b0
   , parameter [4:0]     PF1_BAR1_APERTURE_SIZE=5'b0
   , parameter [4:0]     PF2_BAR1_APERTURE_SIZE=5'b0
   , parameter [4:0]     PF3_BAR1_APERTURE_SIZE=5'b0
   , parameter [2:0]     PF0_BAR2_CONTROL=3'b100
   , parameter [2:0]     PF1_BAR2_CONTROL=3'b100
   , parameter [2:0]     PF2_BAR2_CONTROL=3'b100
   , parameter [2:0]     PF3_BAR2_CONTROL=3'b100
   , parameter [5:0]     PF0_BAR2_APERTURE_SIZE=6'b00011
   , parameter [5:0]     PF1_BAR2_APERTURE_SIZE=6'b00011
   , parameter [5:0]     PF2_BAR2_APERTURE_SIZE=6'b00011
   , parameter [5:0]     PF3_BAR2_APERTURE_SIZE=6'b00011
   , parameter [2:0]     PF0_BAR3_CONTROL=3'b0
   , parameter [2:0]     PF1_BAR3_CONTROL=3'b0
   , parameter [2:0]     PF2_BAR3_CONTROL=3'b0
   , parameter [2:0]     PF3_BAR3_CONTROL=3'b0
   , parameter [4:0]     PF0_BAR3_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF1_BAR3_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF2_BAR3_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF3_BAR3_APERTURE_SIZE=5'b00011
   , parameter [2:0]     PF0_BAR4_CONTROL=3'b100
   , parameter [2:0]     PF1_BAR4_CONTROL=3'b100
   , parameter [2:0]     PF2_BAR4_CONTROL=3'b100
   , parameter [2:0]     PF3_BAR4_CONTROL=3'b100
   , parameter [5:0]     PF0_BAR4_APERTURE_SIZE=6'b00011
   , parameter [5:0]     PF1_BAR4_APERTURE_SIZE=6'b00011
   , parameter [5:0]     PF2_BAR4_APERTURE_SIZE=6'b00011
   , parameter [5:0]     PF3_BAR4_APERTURE_SIZE=6'b00011
   , parameter [2:0]     PF0_BAR5_CONTROL=3'b0
   , parameter [2:0]     PF1_BAR5_CONTROL=3'b0
   , parameter [2:0]     PF2_BAR5_CONTROL=3'b0
   , parameter [2:0]     PF3_BAR5_CONTROL=3'b0
   , parameter [4:0]     PF0_BAR5_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF1_BAR5_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF2_BAR5_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF3_BAR5_APERTURE_SIZE=5'b00011
   , parameter           PF0_EXPANSION_ROM_ENABLE="FALSE"
   , parameter           PF1_EXPANSION_ROM_ENABLE="FALSE"
   , parameter           PF2_EXPANSION_ROM_ENABLE="FALSE"
   , parameter           PF3_EXPANSION_ROM_ENABLE="FALSE"
   , parameter [4:0]     PF0_EXPANSION_ROM_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF1_EXPANSION_ROM_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF2_EXPANSION_ROM_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF3_EXPANSION_ROM_APERTURE_SIZE=5'b00011
   , parameter [7:0]     PF0_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF1_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF2_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF3_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     VFG0_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     VFG1_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     VFG2_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     VFG3_PCIE_CAP_NEXTPTR=8'h0
   , parameter [2:0]     PF0_DEV_CAP_MAX_PAYLOAD_SIZE=3'b011
   , parameter [2:0]     PF1_DEV_CAP_MAX_PAYLOAD_SIZE=3'b011
   , parameter [2:0]     PF2_DEV_CAP_MAX_PAYLOAD_SIZE=3'b011
   , parameter [2:0]     PF3_DEV_CAP_MAX_PAYLOAD_SIZE=3'b011
   , parameter           PF0_DEV_CAP_EXT_TAG_SUPPORTED="TRUE"
   , parameter integer   PF0_DEV_CAP_ENDPOINT_L0S_LATENCY=0
   , parameter integer   PF0_DEV_CAP_ENDPOINT_L1_LATENCY=0
   , parameter           PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE="TRUE"
   , parameter integer   PF0_LINK_CAP_ASPM_SUPPORT=0
   , parameter [0:0]     PF0_LINK_CONTROL_RCB=1'b0
   , parameter           PF0_LINK_STATUS_SLOT_CLOCK_CONFIG="TRUE"
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4=7
   , parameter           PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE="TRUE"
   , parameter           PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT="TRUE"
   , parameter           PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT="TRUE"
   , parameter           PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT="TRUE"
   , parameter           PF0_DEV_CAP2_LTR_SUPPORT="FALSE"
   , parameter           PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT="FALSE"
   , parameter [1:0]     PF0_DEV_CAP2_OBFF_SUPPORT=2'b00
   , parameter           PF0_DEV_CAP2_ARI_FORWARD_ENABLE="FALSE"
   , parameter [7:0]     PF0_MSI_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF1_MSI_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF2_MSI_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF3_MSI_CAP_NEXTPTR=8'h0
   , parameter           PF0_MSI_CAP_PERVECMASKCAP="FALSE"
   , parameter           PF1_MSI_CAP_PERVECMASKCAP="FALSE"
   , parameter           PF2_MSI_CAP_PERVECMASKCAP="FALSE"
   , parameter           PF3_MSI_CAP_PERVECMASKCAP="FALSE"
   , parameter integer   PF0_MSI_CAP_MULTIMSGCAP=0
   , parameter integer   PF1_MSI_CAP_MULTIMSGCAP=0
   , parameter integer   PF2_MSI_CAP_MULTIMSGCAP=0
   , parameter integer   PF3_MSI_CAP_MULTIMSGCAP=0
   , parameter [7:0]     PF0_MSIX_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF1_MSIX_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF2_MSIX_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF3_MSIX_CAP_NEXTPTR=8'h0
   , parameter [7:0]     VFG0_MSIX_CAP_NEXTPTR=PF0_MSIX_CAP_NEXTPTR
   , parameter [7:0]     VFG1_MSIX_CAP_NEXTPTR=PF1_MSIX_CAP_NEXTPTR
   , parameter [7:0]     VFG2_MSIX_CAP_NEXTPTR=PF2_MSIX_CAP_NEXTPTR
   , parameter [7:0]     VFG3_MSIX_CAP_NEXTPTR=PF3_MSIX_CAP_NEXTPTR
   , parameter integer   PF0_MSIX_CAP_PBA_BIR=0
   , parameter integer   PF1_MSIX_CAP_PBA_BIR=0
   , parameter integer   PF2_MSIX_CAP_PBA_BIR=0
   , parameter integer   PF3_MSIX_CAP_PBA_BIR=0
   , parameter integer   VFG0_MSIX_CAP_PBA_BIR=PF0_MSIX_CAP_PBA_BIR
   , parameter integer   VFG1_MSIX_CAP_PBA_BIR=PF1_MSIX_CAP_PBA_BIR
   , parameter integer   VFG2_MSIX_CAP_PBA_BIR=PF2_MSIX_CAP_PBA_BIR
   , parameter integer   VFG3_MSIX_CAP_PBA_BIR=PF3_MSIX_CAP_PBA_BIR
   , parameter [28:0]    PF0_MSIX_CAP_PBA_OFFSET=29'h50
   , parameter [28:0]    PF1_MSIX_CAP_PBA_OFFSET=29'h50
   , parameter [28:0]    PF2_MSIX_CAP_PBA_OFFSET=29'h50
   , parameter [28:0]    PF3_MSIX_CAP_PBA_OFFSET=29'h50
   , parameter [28:0]    VFG0_MSIX_CAP_PBA_OFFSET=PF0_MSIX_CAP_PBA_OFFSET
   , parameter [28:0]    VFG1_MSIX_CAP_PBA_OFFSET=PF1_MSIX_CAP_PBA_OFFSET
   , parameter [28:0]    VFG2_MSIX_CAP_PBA_OFFSET=PF2_MSIX_CAP_PBA_OFFSET
   , parameter [28:0]    VFG3_MSIX_CAP_PBA_OFFSET=PF3_MSIX_CAP_PBA_OFFSET
   , parameter integer   PF0_MSIX_CAP_TABLE_BIR=0
   , parameter integer   PF1_MSIX_CAP_TABLE_BIR=0
   , parameter integer   PF2_MSIX_CAP_TABLE_BIR=0
   , parameter integer   PF3_MSIX_CAP_TABLE_BIR=0
   , parameter integer   VFG0_MSIX_CAP_TABLE_BIR=PF0_MSIX_CAP_TABLE_BIR
   , parameter integer   VFG1_MSIX_CAP_TABLE_BIR=PF1_MSIX_CAP_TABLE_BIR
   , parameter integer   VFG2_MSIX_CAP_TABLE_BIR=PF2_MSIX_CAP_TABLE_BIR
   , parameter integer   VFG3_MSIX_CAP_TABLE_BIR=PF3_MSIX_CAP_TABLE_BIR
   , parameter [28:0]    PF0_MSIX_CAP_TABLE_OFFSET=29'h40
   , parameter [28:0]    PF1_MSIX_CAP_TABLE_OFFSET=29'h40
   , parameter [28:0]    PF2_MSIX_CAP_TABLE_OFFSET=29'h40
   , parameter [28:0]    PF3_MSIX_CAP_TABLE_OFFSET=29'h40
   , parameter [28:0]    VFG0_MSIX_CAP_TABLE_OFFSET=PF0_MSIX_CAP_TABLE_OFFSET
   , parameter [28:0]    VFG1_MSIX_CAP_TABLE_OFFSET=PF1_MSIX_CAP_TABLE_OFFSET
   , parameter [28:0]    VFG2_MSIX_CAP_TABLE_OFFSET=PF2_MSIX_CAP_TABLE_OFFSET
   , parameter [28:0]    VFG3_MSIX_CAP_TABLE_OFFSET=PF3_MSIX_CAP_TABLE_OFFSET
   , parameter [10:0]    PF0_MSIX_CAP_TABLE_SIZE=11'h0
   , parameter [10:0]    PF1_MSIX_CAP_TABLE_SIZE=11'h0
   , parameter [10:0]    PF2_MSIX_CAP_TABLE_SIZE=11'h0
   , parameter [10:0]    PF3_MSIX_CAP_TABLE_SIZE=11'h0
   , parameter [10:0]    VFG0_MSIX_CAP_TABLE_SIZE=PF0_MSIX_CAP_TABLE_SIZE
   , parameter [10:0]    VFG1_MSIX_CAP_TABLE_SIZE=PF1_MSIX_CAP_TABLE_SIZE
   , parameter [10:0]    VFG2_MSIX_CAP_TABLE_SIZE=PF2_MSIX_CAP_TABLE_SIZE
   , parameter [10:0]    VFG3_MSIX_CAP_TABLE_SIZE=PF3_MSIX_CAP_TABLE_SIZE
   , parameter [5:0]     PF0_MSIX_VECTOR_COUNT=6'h4
   , parameter [7:0]     PF0_PM_CAP_ID=8'h1
   , parameter [7:0]     PF0_PM_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF1_PM_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF2_PM_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF3_PM_CAP_NEXTPTR=8'h0
   , parameter           PF0_PM_CAP_PMESUPPORT_D3HOT="TRUE"
   , parameter           PF0_PM_CAP_PMESUPPORT_D1="TRUE"
   , parameter           PF0_PM_CAP_PMESUPPORT_D0="TRUE"
   , parameter           PF0_PM_CAP_SUPP_D1_STATE="TRUE"
   , parameter [2:0]     PF0_PM_CAP_VER_ID=3'h3
   , parameter           PF0_PM_CSR_NOSOFTRESET="TRUE"
   , parameter           PM_ENABLE_L23_ENTRY="TRUE"
   , parameter [7:0]     DNSTREAM_LINK_NUM=8'h0
   , parameter           AUTO_FLR_RESPONSE="FALSE"
   , parameter [11:0]    PF0_DSN_CAP_NEXTPTR=12'h10C
   , parameter [11:0]    PF1_DSN_CAP_NEXTPTR=12'h10C
   , parameter [11:0]    PF2_DSN_CAP_NEXTPTR=12'h10C
   , parameter [11:0]    PF3_DSN_CAP_NEXTPTR=12'h10C
   , parameter           DSN_CAP_ENABLE="FALSE"
   , parameter [3:0]     PF0_VC_CAP_VER=4'h1
   , parameter [11:0]    PF0_VC_CAP_NEXTPTR=12'h0
   , parameter           PF0_VC_CAP_ENABLE="FALSE"
   , parameter [11:0]    PF0_SECONDARY_PCIE_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF0_AER_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF1_AER_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF2_AER_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF3_AER_CAP_NEXTPTR=12'h0
   , parameter           PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE="FALSE"
   , parameter           ARI_CAP_ENABLE="FALSE"
   , parameter [11:0]    PF0_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF1_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF2_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF3_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG0_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG1_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG2_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG3_ARI_CAP_NEXTPTR=12'h0
   , parameter [3:0]     PF0_ARI_CAP_VER=4'h1
   , parameter [7:0]     PF0_ARI_CAP_NEXT_FUNC=8'h0
   , parameter [7:0]     PF1_ARI_CAP_NEXT_FUNC=8'h0
   , parameter [7:0]     PF2_ARI_CAP_NEXT_FUNC=8'h0
   , parameter [7:0]     PF3_ARI_CAP_NEXT_FUNC=8'h0
   , parameter [11:0]    PF0_LTR_CAP_NEXTPTR=12'h0
   , parameter [3:0]     PF0_LTR_CAP_VER=4'h1
   , parameter [9:0]     PF0_LTR_CAP_MAX_SNOOP_LAT=10'h0
   , parameter [9:0]     PF0_LTR_CAP_MAX_NOSNOOP_LAT=10'h0
   , parameter           LTR_TX_MESSAGE_ON_LTR_ENABLE="FALSE"
   , parameter           LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE="FALSE"
   , parameter [9:0]     LTR_TX_MESSAGE_MINIMUM_INTERVAL=10'h250
   , parameter [3:0]     SRIOV_CAP_ENABLE=4'h0
   , parameter [11:0]    PF0_SRIOV_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF1_SRIOV_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF2_SRIOV_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF3_SRIOV_CAP_NEXTPTR=12'h0
   , parameter [3:0]     PF0_SRIOV_CAP_VER=4'h1
   , parameter [3:0]     PF1_SRIOV_CAP_VER=4'h1
   , parameter [3:0]     PF2_SRIOV_CAP_VER=4'h1
   , parameter [3:0]     PF3_SRIOV_CAP_VER=4'h1
   , parameter           PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED="FALSE"
   , parameter           PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED="FALSE"
   , parameter           PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED="FALSE"
   , parameter           PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED="FALSE"
   , parameter [15:0]    PF0_SRIOV_CAP_INITIAL_VF=16'h0
   , parameter [15:0]    PF1_SRIOV_CAP_INITIAL_VF=16'h0
   , parameter [15:0]    PF2_SRIOV_CAP_INITIAL_VF=16'h0
   , parameter [15:0]    PF3_SRIOV_CAP_INITIAL_VF=16'h0
   , parameter [15:0]    PF0_SRIOV_CAP_TOTAL_VF=16'h0
   , parameter [15:0]    PF1_SRIOV_CAP_TOTAL_VF=16'h0
   , parameter [15:0]    PF2_SRIOV_CAP_TOTAL_VF=16'h0
   , parameter [15:0]    PF3_SRIOV_CAP_TOTAL_VF=16'h0
   , parameter [15:0]    PF0_SRIOV_FUNC_DEP_LINK=16'h0
   , parameter [15:0]    PF1_SRIOV_FUNC_DEP_LINK=16'h0
   , parameter [15:0]    PF2_SRIOV_FUNC_DEP_LINK=16'h0
   , parameter [15:0]    PF3_SRIOV_FUNC_DEP_LINK=16'h0
   , parameter [15:0]    PF0_SRIOV_FIRST_VF_OFFSET=16'h0
   , parameter [15:0]    PF1_SRIOV_FIRST_VF_OFFSET=16'h0
   , parameter [15:0]    PF2_SRIOV_FIRST_VF_OFFSET=16'h0
   , parameter [15:0]    PF3_SRIOV_FIRST_VF_OFFSET=16'h0
   , parameter [15:0]    PF0_SRIOV_VF_DEVICE_ID=16'h0
   , parameter [15:0]    PF1_SRIOV_VF_DEVICE_ID=16'h0
   , parameter [15:0]    PF2_SRIOV_VF_DEVICE_ID=16'h0
   , parameter [15:0]    PF3_SRIOV_VF_DEVICE_ID=16'h0
   , parameter [31:0]    PF0_SRIOV_SUPPORTED_PAGE_SIZE=32'h0
   , parameter [31:0]    PF1_SRIOV_SUPPORTED_PAGE_SIZE=32'h0
   , parameter [31:0]    PF2_SRIOV_SUPPORTED_PAGE_SIZE=32'h0
   , parameter [31:0]    PF3_SRIOV_SUPPORTED_PAGE_SIZE=32'h0
   , parameter [2:0]     PF0_SRIOV_BAR0_CONTROL=3'b100
   , parameter [2:0]     PF1_SRIOV_BAR0_CONTROL=3'b100
   , parameter [2:0]     PF2_SRIOV_BAR0_CONTROL=3'b100
   , parameter [2:0]     PF3_SRIOV_BAR0_CONTROL=3'b100
   , parameter [5:0]     PF0_SRIOV_BAR0_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF1_SRIOV_BAR0_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF2_SRIOV_BAR0_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF3_SRIOV_BAR0_APERTURE_SIZE=6'b000011
   , parameter [2:0]     PF0_SRIOV_BAR1_CONTROL=3'b0
   , parameter [2:0]     PF1_SRIOV_BAR1_CONTROL=3'b0
   , parameter [2:0]     PF2_SRIOV_BAR1_CONTROL=3'b0
   , parameter [2:0]     PF3_SRIOV_BAR1_CONTROL=3'b0
   , parameter [4:0]     PF0_SRIOV_BAR1_APERTURE_SIZE=5'b0
   , parameter [4:0]     PF1_SRIOV_BAR1_APERTURE_SIZE=5'b0
   , parameter [4:0]     PF2_SRIOV_BAR1_APERTURE_SIZE=5'b0
   , parameter [4:0]     PF3_SRIOV_BAR1_APERTURE_SIZE=5'b0
   , parameter [2:0]     PF0_SRIOV_BAR2_CONTROL=3'b100
   , parameter [2:0]     PF1_SRIOV_BAR2_CONTROL=3'b100
   , parameter [2:0]     PF2_SRIOV_BAR2_CONTROL=3'b100
   , parameter [2:0]     PF3_SRIOV_BAR2_CONTROL=3'b100
   , parameter [5:0]     PF0_SRIOV_BAR2_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF1_SRIOV_BAR2_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF2_SRIOV_BAR2_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF3_SRIOV_BAR2_APERTURE_SIZE=6'b000011
   , parameter [2:0]     PF0_SRIOV_BAR3_CONTROL=3'b0
   , parameter [2:0]     PF1_SRIOV_BAR3_CONTROL=3'b0
   , parameter [2:0]     PF2_SRIOV_BAR3_CONTROL=3'b0
   , parameter [2:0]     PF3_SRIOV_BAR3_CONTROL=3'b0
   , parameter [4:0]     PF0_SRIOV_BAR3_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF1_SRIOV_BAR3_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF2_SRIOV_BAR3_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF3_SRIOV_BAR3_APERTURE_SIZE=5'b00011
   , parameter [2:0]     PF0_SRIOV_BAR4_CONTROL=3'b100
   , parameter [2:0]     PF1_SRIOV_BAR4_CONTROL=3'b100
   , parameter [2:0]     PF2_SRIOV_BAR4_CONTROL=3'b100
   , parameter [2:0]     PF3_SRIOV_BAR4_CONTROL=3'b100
   , parameter [5:0]     PF0_SRIOV_BAR4_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF1_SRIOV_BAR4_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF2_SRIOV_BAR4_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF3_SRIOV_BAR4_APERTURE_SIZE=6'b000011
   , parameter [2:0]     PF0_SRIOV_BAR5_CONTROL=3'b0
   , parameter [2:0]     PF1_SRIOV_BAR5_CONTROL=3'b0
   , parameter [2:0]     PF2_SRIOV_BAR5_CONTROL=3'b0
   , parameter [2:0]     PF3_SRIOV_BAR5_CONTROL=3'b0
   , parameter [4:0]     PF0_SRIOV_BAR5_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF1_SRIOV_BAR5_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF2_SRIOV_BAR5_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF3_SRIOV_BAR5_APERTURE_SIZE=5'b00011
   , parameter [11:0]    PF0_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF1_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF2_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF3_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG0_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG1_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG2_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG3_TPHR_CAP_NEXTPTR=12'h0
   , parameter [3:0]     PF0_TPHR_CAP_VER=4'h1
   , parameter           PF0_TPHR_CAP_INT_VEC_MODE="TRUE"
   , parameter           PF0_TPHR_CAP_DEV_SPECIFIC_MODE="TRUE"
   , parameter [1:0]     PF0_TPHR_CAP_ST_TABLE_LOC=2'h0
   , parameter [10:0]    PF0_TPHR_CAP_ST_TABLE_SIZE=11'h0
   , parameter [2:0]     PF0_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     PF1_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     PF2_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     PF3_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     VFG0_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     VFG1_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     VFG2_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     VFG3_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter           PF0_TPHR_CAP_ENABLE="FALSE"
   , parameter           TPH_TO_RAM_PIPELINE="TRUE"
   , parameter           TPH_FROM_RAM_PIPELINE="TRUE"
   , parameter           MCAP_ENABLE="FALSE"
   , parameter           MCAP_CONFIGURE_OVERRIDE="FALSE"
   , parameter [11:0]    MCAP_CAP_NEXTPTR=12'h0
   , parameter [15:0]    MCAP_VSEC_ID=16'h0
   , parameter [3:0]     MCAP_VSEC_REV=4'h0
   , parameter [11:0]    MCAP_VSEC_LEN=12'h2C
   , parameter [31:0]    MCAP_FPGA_BITSTREAM_VERSION=32'h0
   , parameter           MCAP_INTERRUPT_ON_MCAP_EOS="FALSE"
   , parameter           MCAP_INTERRUPT_ON_MCAP_ERROR="FALSE"
   , parameter           MCAP_INPUT_GATE_DESIGN_SWITCH="FALSE"
   , parameter           MCAP_EOS_DESIGN_SWITCH="FALSE"
   , parameter           MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH="FALSE"
   , parameter           MCAP_GATE_IO_ENABLE_DESIGN_SWITCH="FALSE"
   , parameter [31:0]    SIM_JTAG_IDCODE=32'h0
   , parameter [7:0]     DEBUG_AXIST_DISABLE_FEATURE_BIT=8'h0
   , parameter           DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS="FALSE"
   , parameter           DEBUG_TL_DISABLE_FC_TIMEOUT="FALSE"
   , parameter           DEBUG_PL_DISABLE_SCRAMBLING="FALSE"
   , parameter           DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL ="FALSE"
   , parameter           DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW ="FALSE"
   , parameter           DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR="FALSE"
   , parameter           DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR="FALSE"
   , parameter           DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR="FALSE"
   , parameter           DEBUG_PL_SIM_RESET_LFSR="FALSE"
   , parameter [15:0]    DEBUG_PL_SPARE=16'h0
   , parameter [15:0]    DEBUG_LL_SPARE=16'h0
   , parameter [15:0]    DEBUG_TL_SPARE=16'h0
   , parameter [15:0]    DEBUG_AXI4ST_SPARE=16'h0
   , parameter [15:0]    DEBUG_CFG_SPARE=16'h0
   , parameter [3:0]     DEBUG_CAR_SPARE=4'h0
   , parameter           TEST_MODE_PIN_CHAR="FALSE"
   , parameter           SPARE_BIT0="FALSE"
   , parameter           SPARE_BIT1=1'b0
   , parameter           SPARE_BIT2=1'b0
   , parameter           SPARE_BIT3="FALSE"
   , parameter           SPARE_BIT4=1'b0
   , parameter           SPARE_BIT5=1'b0
   , parameter           SPARE_BIT6=1'b0
   , parameter           SPARE_BIT7=1'b0
   , parameter           SPARE_BIT8=1'b0
   , parameter [7:0]     SPARE_BYTE0=8'h0
   , parameter [7:0]     SPARE_BYTE1=8'h0
   , parameter [7:0]     SPARE_BYTE2=8'h0
   , parameter [7:0]     SPARE_BYTE3=8'h0
   , parameter [31:0]    SPARE_WORD0=32'h0
   , parameter [31:0]    SPARE_WORD1=32'h0
   , parameter [31:0]    SPARE_WORD2=32'h0
   , parameter [31:0]    SPARE_WORD3=32'h0
   , parameter EXT_PIPE_SIM = "FALSE"

   , parameter PF0_VENDOR_ID='H10EE
   , parameter PF0_SUBSYSTEM_VENDOR_ID='H10EE
   , parameter PF0_DEVICE_ID='H903F
   , parameter PF1_DEVICE_ID='H903F
   , parameter PF2_DEVICE_ID='H903F
   , parameter PF3_DEVICE_ID='H903F
   , parameter PF0_REVISION_ID='H00
   , parameter PF1_REVISION_ID='H00
   , parameter PF2_REVISION_ID='H00
   , parameter PF3_REVISION_ID='H00
   , parameter PF0_SUBSYSTEM_ID='H0007
   , parameter PF1_SUBSYSTEM_ID='H0007
   , parameter PF2_SUBSYSTEM_ID='H0007
   , parameter PF3_SUBSYSTEM_ID='H0007

/// ----------------------------------------------
  , parameter TL_LEGACY_MODE_ENABLE="FALSE",
    parameter DEDICATE_PERST="TRUE",
    parameter SYS_RESET_POLARITY=0,
    parameter DIS_GT_WIZARD="TRUE",
    parameter BMD_PIO_MODE="FALSE",
    parameter COMPLETER_MODEL="FALSE",
    parameter SRIOV_EXD_MODE="FALSE",
    parameter TWO_PORT_SWITCH="FALSE",
    parameter TWO_PORT_CONFIG="X8G3",
    parameter silicon_revision="ES1",
    parameter DEV_PORT_TYPE= 0,
    parameter pcie_blk_locn=0,
    parameter gen_x0y0_xdc=0,
    parameter gen_x0y1_xdc=0,
    parameter gen_x0y2_xdc=0,
    parameter gen_x0y3_xdc=0,
    parameter gen_x0y4_xdc=0,
    parameter gen_x0y5_xdc=0,
    parameter gen_x1y0_xdc=1,
    parameter gen_x1y1_xdc=0,
    parameter gen_x1y2_xdc=0,
    parameter gen_x1y3_xdc=0,
    parameter gen_x1y4_xdc=0,
    parameter gen_x1y5_xdc=0,
    parameter xlnx_ref_board=0,
    parameter PIPE_SIM="FALSE",
    parameter PCIE_FAST_CONFIG="NONE",
    parameter EXT_STARTUP_PRIMITIVE="FALSE",
    parameter PL_INTERFACE="FALSE",
    parameter PCIE_CONFIGURATION="FALSE",
    parameter CFG_STATUS_IF="TRUE",
    parameter TX_FC_IF="TRUE",
    parameter CFG_EXT_IF="TRUE",
    parameter CFG_FC_IF="TRUE",
    parameter PER_FUNC_STATUS_IF="TRUE",
    parameter CFG_MGMT_IF="TRUE",
    parameter CFG_PM_IF="TRUE",
    parameter RCV_MSG_IF="TRUE",
    parameter CFG_TX_MSG_IF="TRUE",
    parameter CFG_CTL_IF="TRUE",
    parameter PCIE_ID_IF="FALSE",
    parameter MSI_EN="TRUE",
    parameter MSIX_EN="FALSE",
    parameter PCIE3_DRP="FALSE",
    parameter TRANSCEIVER_CTRL_STATUS_PORTS="FALSE",
    parameter SHARED_LOGIC=1,
    parameter MCAP_ENABLEMENT="NONE",
    parameter EXT_CH_GT_DRP="FALSE",
    parameter EN_GT_SELECTION="FALSE",
    parameter PLL_TYPE = 0,
    parameter EN_PARITY = "FALSE",
    parameter INS_LOSS_PROFILE = "TRUE",
    parameter MSI_X_OPTIONS="MSI-X_Ext",
    parameter SELECT_QUAD="GTY_Quad_124"
/// ----------------------------------------------

   ) (

    input  wire           pl_gen2_upstream_prefer_deemph
   ,output wire           pl_eq_in_progress
   ,output wire [1:0]     pl_eq_phase
   ,input  wire           pl_redo_eq
   ,input  wire           pl_redo_eq_speed
   ,output wire           pl_eq_mismatch
   ,output wire           pl_redo_eq_pending

   ,output wire [AXI4_DATA_WIDTH-1:0] m_axis_cq_tdata
   ,input  wire [AXI4_DATA_WIDTH-1:0] s_axis_cc_tdata
   ,input  wire [AXI4_DATA_WIDTH-1:0] s_axis_rq_tdata
   ,output wire [AXI4_DATA_WIDTH-1:0] m_axis_rc_tdata
   ,output wire [AXI4_CQ_TUSER_WIDTH-1:0] m_axis_cq_tuser
   ,input  wire [AXI4_CC_TUSER_WIDTH-1:0] s_axis_cc_tuser
   ,output wire           m_axis_cq_tlast
   ,input  wire           s_axis_rq_tlast
   ,output wire           m_axis_rc_tlast
   ,input  wire           s_axis_cc_tlast
   ,input  wire [1:0]     pcie_cq_np_req
   ,output wire [5:0]     pcie_cq_np_req_count
   ,input  wire [AXI4_RQ_TUSER_WIDTH-1:0] s_axis_rq_tuser
   ,output wire [AXI4_RC_TUSER_WIDTH-1:0] m_axis_rc_tuser
   ,output wire [AXI4_TKEEP_WIDTH-1:0] m_axis_cq_tkeep
   ,input  wire [AXI4_TKEEP_WIDTH-1:0] s_axis_cc_tkeep
   ,input  wire [AXI4_TKEEP_WIDTH-1:0] s_axis_rq_tkeep
   ,output wire [AXI4_TKEEP_WIDTH-1:0] m_axis_rc_tkeep
   ,output wire           m_axis_cq_tvalid
   ,input  wire           s_axis_cc_tvalid
   ,input  wire           s_axis_rq_tvalid
   ,output wire           m_axis_rc_tvalid
   ,input  wire           m_axis_cq_tready
   ,output wire [AXI4_CC_TREADY_WIDTH-1:0] s_axis_cc_tready
   ,output wire [AXI4_RQ_TREADY_WIDTH-1:0] s_axis_rq_tready
   ,input  wire           m_axis_rc_tready
   ,output wire [5:0]     pcie_rq_seq_num0
   ,output wire           pcie_rq_seq_num_vld0
   ,output wire [5:0]     pcie_rq_seq_num1
   ,output wire           pcie_rq_seq_num_vld1
   ,output wire [7:0]     pcie_rq_tag0
   ,output wire           pcie_rq_tag_vld0
   ,output wire [7:0]     pcie_rq_tag1
   ,output wire           pcie_rq_tag_vld1
   ,output wire [3:0]     pcie_tfc_nph_av
   ,output wire [3:0]     pcie_tfc_npd_av
   ,output wire [3:0]     pcie_rq_tag_av
   ,input  wire [9:0]     cfg_mgmt_addr
   ,input  wire [7:0]     cfg_mgmt_function_number
   ,input  wire           cfg_mgmt_write
   ,input  wire [31:0]    cfg_mgmt_write_data
   ,input  wire [3:0]     cfg_mgmt_byte_enable
   ,input  wire           cfg_mgmt_read
   ,output wire [31:0]    cfg_mgmt_read_data
   ,output wire           cfg_mgmt_read_write_done
   ,input  wire           cfg_mgmt_debug_access
   ,output wire           cfg_phy_link_down
   ,output wire [1:0]     cfg_phy_link_status
   ,output wire [2:0]     cfg_negotiated_width
   ,output wire [1:0]     cfg_current_speed
   ,output wire [1:0]     cfg_max_payload
   ,output wire [2:0]     cfg_max_read_req
   ,output wire [15:0]    cfg_function_status
   ,output wire [11:0]    cfg_function_power_state
   ,output wire [1:0]     cfg_link_power_state
   ,output wire           cfg_err_cor_out
   ,output wire           cfg_err_nonfatal_out
   ,output wire           cfg_err_fatal_out
   ,output wire           cfg_local_error_valid
   ,output wire [4:0]     cfg_local_error_out
   ,output wire [5:0]     cfg_ltssm_state
   ,output wire [1:0]     cfg_rx_pm_state
   ,output wire [1:0]     cfg_tx_pm_state
   ,output wire [3:0]     cfg_rcb_status
   ,output wire [1:0]     cfg_obff_enable
   ,output wire           cfg_pl_status_change
   ,output wire [3:0]     cfg_tph_requester_enable
   ,output wire [11:0]    cfg_tph_st_mode
   ,output wire           cfg_msg_received
   ,output wire [7:0]     cfg_msg_received_data
   ,output wire [4:0]     cfg_msg_received_type
   ,input  wire           cfg_msg_transmit
   ,input  wire [2:0]     cfg_msg_transmit_type
   ,input  wire [31:0]    cfg_msg_transmit_data
   ,output wire           cfg_msg_transmit_done
   ,output wire [7:0]     cfg_fc_ph
   ,output wire [11:0]    cfg_fc_pd
   ,output wire [7:0]     cfg_fc_nph
   ,output wire [11:0]    cfg_fc_npd
   ,output wire [7:0]     cfg_fc_cplh
   ,output wire [11:0]    cfg_fc_cpld
   ,input  wire [2:0]     cfg_fc_sel
   ,input  wire           cfg_hot_reset_in
   ,output wire           cfg_hot_reset_out
   ,input  wire           cfg_config_space_enable
   ,input  wire [63:0]    cfg_dsn
   ,input  wire [15:0]    cfg_dev_id_pf0
   ,input  wire [15:0]    cfg_dev_id_pf1
   ,input  wire [15:0]    cfg_dev_id_pf2
   ,input  wire [15:0]    cfg_dev_id_pf3
   ,input  wire [15:0]    cfg_vend_id
   ,input  wire [7:0]     cfg_rev_id_pf0
   ,input  wire [7:0]     cfg_rev_id_pf1
   ,input  wire [7:0]     cfg_rev_id_pf2
   ,input  wire [7:0]     cfg_rev_id_pf3
   ,input  wire [15:0]    cfg_subsys_id_pf0
   ,input  wire [15:0]    cfg_subsys_id_pf1
   ,input  wire [15:0]    cfg_subsys_id_pf2
   ,input  wire [15:0]    cfg_subsys_id_pf3
   ,input  wire [15:0]    cfg_subsys_vend_id
   ,input  wire [7:0]     cfg_ds_port_number
   ,input  wire [7:0]     cfg_ds_bus_number
   ,input  wire [4:0]     cfg_ds_device_number
   ,output wire [7:0]     cfg_bus_number
   ,input  wire           cfg_power_state_change_ack
   ,output wire           cfg_power_state_change_interrupt
   ,input  wire           cfg_err_cor_in
   ,input  wire           cfg_err_uncor_in
   ,input  wire [3:0]     cfg_flr_done
   ,output wire [3:0]     cfg_flr_in_process
   ,input  wire           cfg_req_pm_transition_l23_ready
   ,input  wire           cfg_link_training_enable
   ,input  wire [3:0]     cfg_interrupt_int
   ,output wire           cfg_interrupt_sent
   ,input  wire [3:0]     cfg_interrupt_pending
   ,output wire [3:0]     cfg_interrupt_msi_enable
   ,input  wire [31:0]    cfg_interrupt_msi_int
   ,output wire           cfg_interrupt_msi_sent
   ,output wire           cfg_interrupt_msi_fail
   ,output wire [11:0]    cfg_interrupt_msi_mmenable
   ,input  wire [31:0]    cfg_interrupt_msi_pending_status
   ,input  wire [1:0]     cfg_interrupt_msi_pending_status_function_num
   ,input  wire           cfg_interrupt_msi_pending_status_data_enable
   ,output wire           cfg_interrupt_msi_mask_update
   ,input  wire [1:0]     cfg_interrupt_msi_select
   ,output wire [31:0]    cfg_interrupt_msi_data
   ,output wire [3:0]     cfg_interrupt_msix_enable
   ,output wire [3:0]     cfg_interrupt_msix_mask
   ,input  wire [63:0]    cfg_interrupt_msix_address
   ,input  wire [31:0]    cfg_interrupt_msix_data
   ,input  wire           cfg_interrupt_msix_int
   ,input  wire [1:0]     cfg_interrupt_msix_vec_pending
   ,output wire           cfg_interrupt_msix_vec_pending_status
   ,input  wire [2:0]     cfg_interrupt_msi_attr
   ,input  wire           cfg_interrupt_msi_tph_present
   ,input  wire [1:0]     cfg_interrupt_msi_tph_type
   ,input  wire [7:0]     cfg_interrupt_msi_tph_st_tag
   ,input  wire [7:0]     cfg_interrupt_msi_function_number
   ,output wire           cfg_ext_read_received
   ,output wire           cfg_ext_write_received
   ,output wire [9:0]     cfg_ext_register_number
   ,output wire [7:0]     cfg_ext_function_number
   ,output wire [31:0]    cfg_ext_write_data
   ,output wire [3:0]     cfg_ext_write_byte_enable
   ,input  wire [31:0]    cfg_ext_read_data
   ,input  wire           cfg_ext_read_data_valid
   ,output wire [251:0]   cfg_vf_flr_in_process 
   ,input  wire [7:0]     cfg_vf_flr_func_num
   ,input  wire           cfg_vf_flr_done
   ,output wire [503:0]   cfg_vf_status
   ,output wire [755:0]   cfg_vf_power_state
   ,output wire [251:0]   cfg_vf_tph_requester_enable
   ,output wire [755:0]   cfg_vf_tph_st_mode
   ,output wire [251:0]   cfg_interrupt_msix_vf_enable
   ,output wire [251:0]   cfg_interrupt_msix_vf_mask
   ,input  wire           cfg_pm_aspm_l1_entry_reject
   ,input  wire           cfg_pm_aspm_tx_l0s_entry_disable
   ,input  wire [1:0]     conf_req_type
   ,input  wire [3:0]     conf_req_reg_num
   ,input  wire [31:0]    conf_req_data
   ,input  wire           conf_req_valid
   ,output wire           conf_req_ready
   ,output wire [31:0]    conf_resp_rdata
   ,output wire           conf_resp_valid
   ,output wire           conf_mcap_design_switch
   ,output wire           conf_mcap_eos
   ,output wire           conf_mcap_in_use_by_pcie
   ,input  wire           conf_mcap_request_by_conf
   ,output wire           user_clk
   ,output wire           user_reset
   ,output wire           user_lnk_up
   ,input  wire           sys_clk
   ,input  wire           sys_clk_gt
   ,input  wire           sys_reset
   ,input  wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]     pci_exp_rxp
   ,input  wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]     pci_exp_rxn
   ,output wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]     pci_exp_txp
   ,output wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]     pci_exp_txn
  // PIPE INTERFACE
   ,input  wire  [25:0] common_commands_in
   ,input  wire [83:0]  pipe_rx_0_sigs
   ,input  wire [83:0]  pipe_rx_1_sigs
   ,input  wire [83:0]  pipe_rx_2_sigs
   ,input  wire [83:0]  pipe_rx_3_sigs
   ,input  wire [83:0]  pipe_rx_4_sigs
   ,input  wire [83:0]  pipe_rx_5_sigs
   ,input  wire [83:0]  pipe_rx_6_sigs
   ,input  wire [83:0]  pipe_rx_7_sigs
   ,input  wire [83:0]  pipe_rx_8_sigs
   ,input  wire [83:0]  pipe_rx_9_sigs
   ,input  wire [83:0]  pipe_rx_10_sigs
   ,input  wire [83:0]  pipe_rx_11_sigs
   ,input  wire [83:0]  pipe_rx_12_sigs
   ,input  wire [83:0]  pipe_rx_13_sigs
   ,input  wire [83:0]  pipe_rx_14_sigs
   ,input  wire [83:0]  pipe_rx_15_sigs
                      
   ,output wire [16:0]  common_commands_out
   ,output wire [69:0]  pipe_tx_0_sigs
   ,output wire [69:0]  pipe_tx_1_sigs
   ,output wire [69:0]  pipe_tx_2_sigs
   ,output wire [69:0]  pipe_tx_3_sigs
   ,output wire [69:0]  pipe_tx_4_sigs
   ,output wire [69:0]  pipe_tx_5_sigs
   ,output wire [69:0]  pipe_tx_6_sigs
   ,output wire [69:0]  pipe_tx_7_sigs
   ,output  wire [69:0]  pipe_tx_8_sigs
   ,output  wire [69:0]  pipe_tx_9_sigs
   ,output  wire [69:0]  pipe_tx_10_sigs
   ,output  wire [69:0]  pipe_tx_11_sigs
   ,output  wire [69:0]  pipe_tx_12_sigs
   ,output  wire [69:0]  pipe_tx_13_sigs
   ,output  wire [69:0]  pipe_tx_14_sigs
   ,output  wire [69:0]  pipe_tx_15_sigs
  );

   wire           pcie_perst0_b;
   wire           pcie_perst1_b;
   wire           sys_clk_bufg;
   wire           phy_rdy ;
   wire           phy_rdy_phystatus;
   wire [1:0]     pipe_rx00_char_is_k;
   wire [1:0]     pipe_rx01_char_is_k;
   wire [1:0]     pipe_rx02_char_is_k;
   wire [1:0]     pipe_rx03_char_is_k;
   wire [1:0]     pipe_rx04_char_is_k;
   wire [1:0]     pipe_rx05_char_is_k;
   wire [1:0]     pipe_rx06_char_is_k;
   wire [1:0]     pipe_rx07_char_is_k;
   wire [1:0]     pipe_rx08_char_is_k;
   wire [1:0]     pipe_rx09_char_is_k;
   wire [1:0]     pipe_rx10_char_is_k;
   wire [1:0]     pipe_rx11_char_is_k;
   wire [1:0]     pipe_rx12_char_is_k;
   wire [1:0]     pipe_rx13_char_is_k;
   wire [1:0]     pipe_rx14_char_is_k;
   wire [1:0]     pipe_rx15_char_is_k;
   wire           pipe_rx00_valid;
   wire           pipe_rx01_valid;
   wire           pipe_rx02_valid;
   wire           pipe_rx03_valid;
   wire           pipe_rx04_valid;
   wire           pipe_rx05_valid;
   wire           pipe_rx06_valid;
   wire           pipe_rx07_valid;
   wire           pipe_rx08_valid;
   wire           pipe_rx09_valid;
   wire           pipe_rx10_valid;
   wire           pipe_rx11_valid;
   wire           pipe_rx12_valid;
   wire           pipe_rx13_valid;
   wire           pipe_rx14_valid;
   wire           pipe_rx15_valid;
   wire [63:0]    pipe_rx00_data;
   wire [63:0]    pipe_rx01_data;
   wire [63:0]    pipe_rx02_data;
   wire [63:0]    pipe_rx03_data;
   wire [63:0]    pipe_rx04_data;
   wire [63:0]    pipe_rx05_data;
   wire [63:0]    pipe_rx06_data;
   wire [63:0]    pipe_rx07_data;
   wire [63:0]    pipe_rx08_data;
   wire [63:0]    pipe_rx09_data;
   wire [63:0]    pipe_rx10_data;
   wire [63:0]    pipe_rx11_data;
   wire [63:0]    pipe_rx12_data;
   wire [63:0]    pipe_rx13_data;
   wire [63:0]    pipe_rx14_data;
   wire [63:0]    pipe_rx15_data;
   wire           pipe_rx00_polarity;
   wire           pipe_rx01_polarity;
   wire           pipe_rx02_polarity;
   wire           pipe_rx03_polarity;
   wire           pipe_rx04_polarity;
   wire           pipe_rx05_polarity;
   wire           pipe_rx06_polarity;
   wire           pipe_rx07_polarity;
   wire           pipe_rx08_polarity;
   wire           pipe_rx09_polarity;
   wire           pipe_rx10_polarity;
   wire           pipe_rx11_polarity;
   wire           pipe_rx12_polarity;
   wire           pipe_rx13_polarity;
   wire           pipe_rx14_polarity;
   wire           pipe_rx15_polarity;
   wire [2:0]     pipe_rx00_status;
   wire [2:0]     pipe_rx01_status;
   wire [2:0]     pipe_rx02_status;
   wire [2:0]     pipe_rx03_status;
   wire [2:0]     pipe_rx04_status;
   wire [2:0]     pipe_rx05_status;
   wire [2:0]     pipe_rx06_status;
   wire [2:0]     pipe_rx07_status;
   wire [2:0]     pipe_rx08_status;
   wire [2:0]     pipe_rx09_status;
   wire [2:0]     pipe_rx10_status;
   wire [2:0]     pipe_rx11_status;
   wire [2:0]     pipe_rx12_status;
   wire [2:0]     pipe_rx13_status;
   wire [2:0]     pipe_rx14_status;
   wire [2:0]     pipe_rx15_status;
   wire           pipe_rx00_phy_status;
   wire           pipe_rx01_phy_status;
   wire           pipe_rx02_phy_status;
   wire           pipe_rx03_phy_status;
   wire           pipe_rx04_phy_status;
   wire           pipe_rx05_phy_status;
   wire           pipe_rx06_phy_status;
   wire           pipe_rx07_phy_status;
   wire           pipe_rx08_phy_status;
   wire           pipe_rx09_phy_status;
   wire           pipe_rx10_phy_status;
   wire           pipe_rx11_phy_status;
   wire           pipe_rx12_phy_status;
   wire           pipe_rx13_phy_status;
   wire           pipe_rx14_phy_status;
   wire           pipe_rx15_phy_status;
   wire           pipe_rx00_elec_idle;
   wire           pipe_rx01_elec_idle;
   wire           pipe_rx02_elec_idle;
   wire           pipe_rx03_elec_idle;
   wire           pipe_rx04_elec_idle;
   wire           pipe_rx05_elec_idle;
   wire           pipe_rx06_elec_idle;
   wire           pipe_rx07_elec_idle;
   wire           pipe_rx08_elec_idle;
   wire           pipe_rx09_elec_idle;
   wire           pipe_rx10_elec_idle;
   wire           pipe_rx11_elec_idle;
   wire           pipe_rx12_elec_idle;
   wire           pipe_rx13_elec_idle;
   wire           pipe_rx14_elec_idle;
   wire           pipe_rx15_elec_idle;
   wire           pipe_rx00_data_valid;
   wire           pipe_rx01_data_valid;
   wire           pipe_rx02_data_valid;
   wire           pipe_rx03_data_valid;
   wire           pipe_rx04_data_valid;
   wire           pipe_rx05_data_valid;
   wire           pipe_rx06_data_valid;
   wire           pipe_rx07_data_valid;
   wire           pipe_rx08_data_valid;
   wire           pipe_rx09_data_valid;
   wire           pipe_rx10_data_valid;
   wire           pipe_rx11_data_valid;
   wire           pipe_rx12_data_valid;
   wire           pipe_rx13_data_valid;
   wire           pipe_rx14_data_valid;
   wire           pipe_rx15_data_valid;
   wire [1:0]     pipe_rx00_start_block;
   wire [1:0]     pipe_rx01_start_block;
   wire [1:0]     pipe_rx02_start_block;
   wire [1:0]     pipe_rx03_start_block;
   wire [1:0]     pipe_rx04_start_block;
   wire [1:0]     pipe_rx05_start_block;
   wire [1:0]     pipe_rx06_start_block;
   wire [1:0]     pipe_rx07_start_block;
   wire [1:0]     pipe_rx08_start_block;
   wire [1:0]     pipe_rx09_start_block;
   wire [1:0]     pipe_rx10_start_block;
   wire [1:0]     pipe_rx11_start_block;
   wire [1:0]     pipe_rx12_start_block;
   wire [1:0]     pipe_rx13_start_block;
   wire [1:0]     pipe_rx14_start_block;
   wire [1:0]     pipe_rx15_start_block;
   wire [1:0]     pipe_rx00_sync_header;
   wire [1:0]     pipe_rx01_sync_header;
   wire [1:0]     pipe_rx02_sync_header;
   wire [1:0]     pipe_rx03_sync_header;
   wire [1:0]     pipe_rx04_sync_header;
   wire [1:0]     pipe_rx05_sync_header;
   wire [1:0]     pipe_rx06_sync_header;
   wire [1:0]     pipe_rx07_sync_header;
   wire [1:0]     pipe_rx08_sync_header;
   wire [1:0]     pipe_rx09_sync_header;
   wire [1:0]     pipe_rx10_sync_header;
   wire [1:0]     pipe_rx11_sync_header;
   wire [1:0]     pipe_rx12_sync_header;
   wire [1:0]     pipe_rx13_sync_header;
   wire [1:0]     pipe_rx14_sync_header;
   wire [1:0]     pipe_rx15_sync_header;
   wire           pipe_tx00_compliance;
   wire           pipe_tx01_compliance;
   wire           pipe_tx02_compliance;
   wire           pipe_tx03_compliance;
   wire           pipe_tx04_compliance;
   wire           pipe_tx05_compliance;
   wire           pipe_tx06_compliance;
   wire           pipe_tx07_compliance;
   wire           pipe_tx08_compliance;
   wire           pipe_tx09_compliance;
   wire           pipe_tx10_compliance;
   wire           pipe_tx11_compliance;
   wire           pipe_tx12_compliance;
   wire           pipe_tx13_compliance;
   wire           pipe_tx14_compliance;
   wire           pipe_tx15_compliance;
   wire [1:0]     pipe_tx00_char_is_k;
   wire [1:0]     pipe_tx01_char_is_k;
   wire [1:0]     pipe_tx02_char_is_k;
   wire [1:0]     pipe_tx03_char_is_k;
   wire [1:0]     pipe_tx04_char_is_k;
   wire [1:0]     pipe_tx05_char_is_k;
   wire [1:0]     pipe_tx06_char_is_k;
   wire [1:0]     pipe_tx07_char_is_k;
   wire [1:0]     pipe_tx08_char_is_k;
   wire [1:0]     pipe_tx09_char_is_k;
   wire [1:0]     pipe_tx10_char_is_k;
   wire [1:0]     pipe_tx11_char_is_k;
   wire [1:0]     pipe_tx12_char_is_k;
   wire [1:0]     pipe_tx13_char_is_k;
   wire [1:0]     pipe_tx14_char_is_k;
   wire [1:0]     pipe_tx15_char_is_k;
   wire [31:0]    pipe_tx00_data;
   wire [31:0]    pipe_tx01_data;
   wire [31:0]    pipe_tx02_data;
   wire [31:0]    pipe_tx03_data;
   wire [31:0]    pipe_tx04_data;
   wire [31:0]    pipe_tx05_data;
   wire [31:0]    pipe_tx06_data;
   wire [31:0]    pipe_tx07_data;
   wire [31:0]    pipe_tx08_data;
   wire [31:0]    pipe_tx09_data;
   wire [31:0]    pipe_tx10_data;
   wire [31:0]    pipe_tx11_data;
   wire [31:0]    pipe_tx12_data;
   wire [31:0]    pipe_tx13_data;
   wire [31:0]    pipe_tx14_data;
   wire [31:0]    pipe_tx15_data;
   wire           pipe_tx00_elec_idle;
   wire           pipe_tx01_elec_idle;
   wire           pipe_tx02_elec_idle;
   wire           pipe_tx03_elec_idle;
   wire           pipe_tx04_elec_idle;
   wire           pipe_tx05_elec_idle;
   wire           pipe_tx06_elec_idle;
   wire           pipe_tx07_elec_idle;
   wire           pipe_tx08_elec_idle;
   wire           pipe_tx09_elec_idle;
   wire           pipe_tx10_elec_idle;
   wire           pipe_tx11_elec_idle;
   wire           pipe_tx12_elec_idle;
   wire           pipe_tx13_elec_idle;
   wire           pipe_tx14_elec_idle;
   wire           pipe_tx15_elec_idle;
   wire [1:0]     pipe_tx00_powerdown;
   wire [1:0]     pipe_tx01_powerdown;
   wire [1:0]     pipe_tx02_powerdown;
   wire [1:0]     pipe_tx03_powerdown;
   wire [1:0]     pipe_tx04_powerdown;
   wire [1:0]     pipe_tx05_powerdown;
   wire [1:0]     pipe_tx06_powerdown;
   wire [1:0]     pipe_tx07_powerdown;
   wire [1:0]     pipe_tx08_powerdown;
   wire [1:0]     pipe_tx09_powerdown;
   wire [1:0]     pipe_tx10_powerdown;
   wire [1:0]     pipe_tx11_powerdown;
   wire [1:0]     pipe_tx12_powerdown;
   wire [1:0]     pipe_tx13_powerdown;
   wire [1:0]     pipe_tx14_powerdown;
   wire [1:0]     pipe_tx15_powerdown;
   wire           pipe_tx00_data_valid;
   wire           pipe_tx01_data_valid;
   wire           pipe_tx02_data_valid;
   wire           pipe_tx03_data_valid;
   wire           pipe_tx04_data_valid;
   wire           pipe_tx05_data_valid;
   wire           pipe_tx06_data_valid;
   wire           pipe_tx07_data_valid;
   wire           pipe_tx08_data_valid;
   wire           pipe_tx09_data_valid;
   wire           pipe_tx10_data_valid;
   wire           pipe_tx11_data_valid;
   wire           pipe_tx12_data_valid;
   wire           pipe_tx13_data_valid;
   wire           pipe_tx14_data_valid;
   wire           pipe_tx15_data_valid;
   wire           pipe_tx00_start_block;
   wire           pipe_tx01_start_block;
   wire           pipe_tx02_start_block;
   wire           pipe_tx03_start_block;
   wire           pipe_tx04_start_block;
   wire           pipe_tx05_start_block;
   wire           pipe_tx06_start_block;
   wire           pipe_tx07_start_block;
   wire           pipe_tx08_start_block;
   wire           pipe_tx09_start_block;
   wire           pipe_tx10_start_block;
   wire           pipe_tx11_start_block;
   wire           pipe_tx12_start_block;
   wire           pipe_tx13_start_block;
   wire           pipe_tx14_start_block;
   wire           pipe_tx15_start_block;
   wire [1:0]     pipe_tx00_sync_header;
   wire [1:0]     pipe_tx01_sync_header;
   wire [1:0]     pipe_tx02_sync_header;
   wire [1:0]     pipe_tx03_sync_header;
   wire [1:0]     pipe_tx04_sync_header;
   wire [1:0]     pipe_tx05_sync_header;
   wire [1:0]     pipe_tx06_sync_header;
   wire [1:0]     pipe_tx07_sync_header;
   wire [1:0]     pipe_tx08_sync_header;
   wire [1:0]     pipe_tx09_sync_header;
   wire [1:0]     pipe_tx10_sync_header;
   wire [1:0]     pipe_tx11_sync_header;
   wire [1:0]     pipe_tx12_sync_header;
   wire [1:0]     pipe_tx13_sync_header;
   wire [1:0]     pipe_tx14_sync_header;
   wire [1:0]     pipe_tx15_sync_header;
   wire [1:0]     pipe_rx00_eq_control;
   wire [1:0]     pipe_rx01_eq_control;
   wire [1:0]     pipe_rx02_eq_control;
   wire [1:0]     pipe_rx03_eq_control;
   wire [1:0]     pipe_rx04_eq_control;
   wire [1:0]     pipe_rx05_eq_control;
   wire [1:0]     pipe_rx06_eq_control;
   wire [1:0]     pipe_rx07_eq_control;
   wire [1:0]     pipe_rx08_eq_control;
   wire [1:0]     pipe_rx09_eq_control;
   wire [1:0]     pipe_rx10_eq_control;
   wire [1:0]     pipe_rx11_eq_control;
   wire [1:0]     pipe_rx12_eq_control;
   wire [1:0]     pipe_rx13_eq_control;
   wire [1:0]     pipe_rx14_eq_control;
   wire [1:0]     pipe_rx15_eq_control;
   wire           pipe_rx00_eq_lp_lf_fs_sel;
   wire           pipe_rx01_eq_lp_lf_fs_sel;
   wire           pipe_rx02_eq_lp_lf_fs_sel;
   wire           pipe_rx03_eq_lp_lf_fs_sel;
   wire           pipe_rx04_eq_lp_lf_fs_sel;
   wire           pipe_rx05_eq_lp_lf_fs_sel;
   wire           pipe_rx06_eq_lp_lf_fs_sel;
   wire           pipe_rx07_eq_lp_lf_fs_sel;
   wire           pipe_rx08_eq_lp_lf_fs_sel;
   wire           pipe_rx09_eq_lp_lf_fs_sel;
   wire           pipe_rx10_eq_lp_lf_fs_sel;
   wire           pipe_rx11_eq_lp_lf_fs_sel;
   wire           pipe_rx12_eq_lp_lf_fs_sel;
   wire           pipe_rx13_eq_lp_lf_fs_sel;
   wire           pipe_rx14_eq_lp_lf_fs_sel;
   wire           pipe_rx15_eq_lp_lf_fs_sel;
   wire [17:0]    pipe_rx00_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx01_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx02_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx03_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx04_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx05_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx06_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx07_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx08_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx09_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx10_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx11_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx12_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx13_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx14_eq_lp_new_tx_coeff_or_preset;
   wire [17:0]    pipe_rx15_eq_lp_new_tx_coeff_or_preset;
   wire           pipe_rx00_eq_lp_adapt_done;
   wire           pipe_rx01_eq_lp_adapt_done;
   wire           pipe_rx02_eq_lp_adapt_done;
   wire           pipe_rx03_eq_lp_adapt_done;
   wire           pipe_rx04_eq_lp_adapt_done;
   wire           pipe_rx05_eq_lp_adapt_done;
   wire           pipe_rx06_eq_lp_adapt_done;
   wire           pipe_rx07_eq_lp_adapt_done;
   wire           pipe_rx08_eq_lp_adapt_done;
   wire           pipe_rx09_eq_lp_adapt_done;
   wire           pipe_rx10_eq_lp_adapt_done;
   wire           pipe_rx11_eq_lp_adapt_done;
   wire           pipe_rx12_eq_lp_adapt_done;
   wire           pipe_rx13_eq_lp_adapt_done;
   wire           pipe_rx14_eq_lp_adapt_done;
   wire           pipe_rx15_eq_lp_adapt_done;
   wire           pipe_rx00_eq_done;
   wire           pipe_rx01_eq_done;
   wire           pipe_rx02_eq_done;
   wire           pipe_rx03_eq_done;
   wire           pipe_rx04_eq_done;
   wire           pipe_rx05_eq_done;
   wire           pipe_rx06_eq_done;
   wire           pipe_rx07_eq_done;
   wire           pipe_rx08_eq_done;
   wire           pipe_rx09_eq_done;
   wire           pipe_rx10_eq_done;
   wire           pipe_rx11_eq_done;
   wire           pipe_rx12_eq_done;
   wire           pipe_rx13_eq_done;
   wire           pipe_rx14_eq_done;
   wire           pipe_rx15_eq_done;
   wire [1:0]     pipe_tx00_eq_control;
   wire [1:0]     pipe_tx01_eq_control;
   wire [1:0]     pipe_tx02_eq_control;
   wire [1:0]     pipe_tx03_eq_control;
   wire [1:0]     pipe_tx04_eq_control;
   wire [1:0]     pipe_tx05_eq_control;
   wire [1:0]     pipe_tx06_eq_control;
   wire [1:0]     pipe_tx07_eq_control;
   wire [1:0]     pipe_tx08_eq_control;
   wire [1:0]     pipe_tx09_eq_control;
   wire [1:0]     pipe_tx10_eq_control;
   wire [1:0]     pipe_tx11_eq_control;
   wire [1:0]     pipe_tx12_eq_control;
   wire [1:0]     pipe_tx13_eq_control;
   wire [1:0]     pipe_tx14_eq_control;
   wire [1:0]     pipe_tx15_eq_control;
   wire [5:0]     pipe_tx00_eq_deemph;
   wire [5:0]     pipe_tx01_eq_deemph;
   wire [5:0]     pipe_tx02_eq_deemph;
   wire [5:0]     pipe_tx03_eq_deemph;
   wire [5:0]     pipe_tx04_eq_deemph;
   wire [5:0]     pipe_tx05_eq_deemph;
   wire [5:0]     pipe_tx06_eq_deemph;
   wire [5:0]     pipe_tx07_eq_deemph;
   wire [5:0]     pipe_tx08_eq_deemph;
   wire [5:0]     pipe_tx09_eq_deemph;
   wire [5:0]     pipe_tx10_eq_deemph;
   wire [5:0]     pipe_tx11_eq_deemph;
   wire [5:0]     pipe_tx12_eq_deemph;
   wire [5:0]     pipe_tx13_eq_deemph;
   wire [5:0]     pipe_tx14_eq_deemph;
   wire [5:0]     pipe_tx15_eq_deemph;
   wire [17:0]    pipe_tx00_eq_coeff;
   wire [17:0]    pipe_tx01_eq_coeff;
   wire [17:0]    pipe_tx02_eq_coeff;
   wire [17:0]    pipe_tx03_eq_coeff;
   wire [17:0]    pipe_tx04_eq_coeff;
   wire [17:0]    pipe_tx05_eq_coeff;
   wire [17:0]    pipe_tx06_eq_coeff;
   wire [17:0]    pipe_tx07_eq_coeff;
   wire [17:0]    pipe_tx08_eq_coeff;
   wire [17:0]    pipe_tx09_eq_coeff;
   wire [17:0]    pipe_tx10_eq_coeff;
   wire [17:0]    pipe_tx11_eq_coeff;
   wire [17:0]    pipe_tx12_eq_coeff;
   wire [17:0]    pipe_tx13_eq_coeff;
   wire [17:0]    pipe_tx14_eq_coeff;
   wire [17:0]    pipe_tx15_eq_coeff;
   wire           pipe_tx00_eq_done;
   wire           pipe_tx01_eq_done;
   wire           pipe_tx02_eq_done;
   wire           pipe_tx03_eq_done;
   wire           pipe_tx04_eq_done;
   wire           pipe_tx05_eq_done;
   wire           pipe_tx06_eq_done;
   wire           pipe_tx07_eq_done;
   wire           pipe_tx08_eq_done;
   wire           pipe_tx09_eq_done;
   wire           pipe_tx10_eq_done;
   wire           pipe_tx11_eq_done;
   wire           pipe_tx12_eq_done;
   wire           pipe_tx13_eq_done;
   wire           pipe_tx14_eq_done;
   wire           pipe_tx15_eq_done;

   wire [3:0]     pipe_rx_eq_lp_tx_preset;
   wire [5:0]     pipe_rx_eq_lp_lf_fs;
   wire           pipe_tx_rcvr_det;
   wire [1:0]     pipe_tx_rate;
   reg  [1:0]     pipe_tx_rate_ff;
   reg            speed_change_in_progress;
   wire           pipe_tx_deemph;
   wire [2:0]     pipe_tx_margin;
   wire           pipe_tx_swing;
   wire           pipe_tx_reset;
   wire [5:0]     pipe_eq_fs;
   wire [5:0]     pipe_eq_lf;

   wire [2:0]     pipe_rx_eq_preset = 3'b0;

   wire           user_clk_en;
   wire           core_clk;
   wire           sys_rst_n;
   wire           sys_or_hot_rst;
   wire           user_lnk_up_int;
   wire           user_clk2 = (AXISTEN_IF_EXT_512 == "TRUE") ? core_clk : user_clk;
   wire           mcap_clk;
   wire		        pipe_clk;   



   wire [(PL_LINK_CAP_MAX_LINK_WIDTH*64)-1:0]     PHY_RXDATA;
   wire [(PL_LINK_CAP_MAX_LINK_WIDTH* 2)-1:0]     PHY_RXDATAK;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          PHY_RXDATA_VALID;
   wire [(PL_LINK_CAP_MAX_LINK_WIDTH* 2)-1:0]     PHY_RXSTART_BLOCK;
   reg [(PL_LINK_CAP_MAX_LINK_WIDTH* 2)-1:0]     PHY_RXSYNC_HEADER;

   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          PHY_RXVALID;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          PHY_PHYSTATUS;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          phy_status_fix;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          PHY_RXELECIDLE;
   wire [(PL_LINK_CAP_MAX_LINK_WIDTH*3)-1:0]      PHY_RXSTATUS;

   wire [(PL_LINK_CAP_MAX_LINK_WIDTH*18)-1:0]     PHY_TXEQ_NEW_COEFF;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          PHY_TXEQ_DONE;

   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          PHY_RXEQ_LFFS_SEL;
   wire [(PL_LINK_CAP_MAX_LINK_WIDTH*18)-1:0]     PHY_RXEQ_NEW_TXCOEFF;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          PHY_RXEQ_ADAPT_DONE;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          PHY_RXEQ_DONE;

   wire [PL_LINK_CAP_MAX_LINK_WIDTH*64-1:0]       PHY_TXDATA;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH*2-1:0]        PHY_TXDATAK;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          PHY_TXDATA_VALID;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          PHY_TXSTART_BLOCK;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH*2-1:0]        PHY_TXSYNC_HEADER;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          PHY_TXELECIDLE;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          PHY_TXCOMPLIANCE;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH-1:0]          PHY_RXPOLARITY;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH*2-1:0]        PHY_TXEQ_CTRL;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH*4-1:0]        PHY_TXEQ_PRESET;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH*6-1:0]        PHY_TXEQ_COEFF;
   wire [PL_LINK_CAP_MAX_LINK_WIDTH*2-1:0]        PHY_RXEQ_CTRL;

(* keep = "true", max_fanout = 800 *) reg   reg_user_lnk_up;
(* keep = "true", max_fanout = 800 *) reg   user_reset_int;
(* keep = "true", max_fanout = 800 *) reg   reg_user_reset;

   reg   as_cdr_hold_req_user;
   reg   as_cdr_hold_req_ff;
   reg   as_cdr_hold_req_ff1;
   reg   as_mac_in_detect_user;
   reg   as_mac_in_detect_ff;
   reg   as_mac_in_detect_ff1;

// Gate rxsync_header with rxstart_block
wire [(PL_LINK_CAP_MAX_LINK_WIDTH* 2)-1:0]     rxsync_header_nogate;
integer ii;
always @*
  for (ii=0;ii<(PL_LINK_CAP_MAX_LINK_WIDTH*2);ii=ii+2)
    PHY_RXSYNC_HEADER[ii+:2] = rxsync_header_nogate[ii+:2] & {2{^PHY_RXSTART_BLOCK[ii+:2]}};


// Workaround for the double-triggering on cfg_msg_transmit
wire cfg_msg_transmit_int = cfg_msg_transmit & ~cfg_msg_transmit_done;

generate if (EXT_PIPE_SIM == "TRUE") 
begin
  /////////////// phy_rdy, rcvr det , seepd_change & gt_powerdown /////////////////////////////
  
  reg [31:0] phy_rdy_reg = 32'b0;
  reg [31:0] rcvr_det_reg     = 32'b0;
  reg  [7:0] pipe_rate_reg    = 8'b0;
  reg  [7:0] gt_powerdown_reg = {4{2'b10}};
  
  wire      rcvr_det;
  wire      speed_change;
  wire      gt_powerdown;

  wire      pipe_tx0_rcvr_det;

    
  always @ (posedge pipe_clk)
  begin
   phy_rdy_reg      <= {phy_rdy_reg[30:0], sys_rst_n};
   rcvr_det_reg     <= {rcvr_det_reg[30:0], pipe_tx0_rcvr_det};
   pipe_rate_reg    <= {pipe_rate_reg[5:0], common_commands_out[2:1]};
   gt_powerdown_reg <= {gt_powerdown_reg[5:0],pipe_tx_0_sigs[41:40]};
  end 
  
  assign phy_rdy      =  phy_rdy_reg[31];
  assign rcvr_det     = ~rcvr_det_reg[30] && rcvr_det_reg[29];
  assign speed_change = (pipe_rate_reg[7:6] != pipe_rate_reg[5:4])? 1'b1 : 1'b0;
  assign gt_powerdown = (gt_powerdown_reg[7:6] == 2'b10 && gt_powerdown_reg[5:4] == 2'b0)? 1'b1 : 1'b0;
  
  
  
  //////// generate Rx status and Phy status ////////////// 
  
  wire [2:0] rx_status;
  wire       phy_status;
  
  assign  rx_status  = (pipe_tx0_rcvr_det && rcvr_det) ? 3'b011 : 3'b0;
  assign  phy_status = (pipe_tx0_rcvr_det && rcvr_det) || speed_change || gt_powerdown ;

   
  //////// generate clocks for pipe mode //////////////
 
  wire clk_500;
  wire clk_250;
  wire clk_125;
  wire clk_62_5;
 
  xp4_usp_smsw_sys_clk_gen_ps 	#(.offset(7000),.halfcycle(1000)) clk_gen_500  (.sys_clk(clk_500));
  xp4_usp_smsw_sys_clk_gen_ps 	#(.offset(6000),.halfcycle(2000)) clk_gen_250  (.sys_clk(clk_250));
  xp4_usp_smsw_sys_clk_gen_ps 	#(.offset(4000),.halfcycle(4000)) clk_gen_125  (.sys_clk(clk_125));
  xp4_usp_smsw_sys_clk_gen_ps 	#(.offset(0000),.halfcycle(8000)) clk_gen_62_5 (.sys_clk(clk_62_5));
 
  assign mcap_clk = (CRM_USER_CLK_FREQ == 2'b10 || CRM_USER_CLK_FREQ == 2'b11) ? clk_125 : user_clk;
  assign pipe_clk = (common_commands_out[2:1] == 2'b0)? clk_125 : clk_250;
  assign core_clk = (CRM_CORE_CLK_FREQ_500 == "TRUE") ? clk_500 : clk_250 ;
  assign user_clk = (CRM_USER_CLK_FREQ == 2'b10 || CRM_USER_CLK_FREQ == 2'b11) ? clk_250: ((CRM_USER_CLK_FREQ == 01) ? clk_125 : clk_62_5);

  // PCIE_4_0 Instance
  xp4_usp_smsw_pipe 
  #(

    .TCQ(TCQ)
   ,.IMPL_TARGET(IMPL_TARGET)
   ,.AXISTEN_IF_EXT_512_INTFC_RAM_STYLE(AXISTEN_IF_EXT_512_INTFC_RAM_STYLE)
   ,.CRM_CORE_CLK_FREQ_500(CRM_CORE_CLK_FREQ_500)
   ,.CRM_USER_CLK_FREQ(CRM_USER_CLK_FREQ)
   ,.AXISTEN_IF_WIDTH(AXISTEN_IF_WIDTH)
   ,.AXISTEN_IF_EXT_512_CQ_STRADDLE(AXISTEN_IF_EXT_512_CQ_STRADDLE)
   ,.AXISTEN_IF_EXT_512_CC_STRADDLE(AXISTEN_IF_EXT_512_CC_STRADDLE)
   ,.AXISTEN_IF_EXT_512_RQ_STRADDLE(AXISTEN_IF_EXT_512_RQ_STRADDLE)
   ,.AXISTEN_IF_EXT_512_RC_STRADDLE(AXISTEN_IF_EXT_512_RC_STRADDLE)
   ,.AXISTEN_IF_EXT_512_RC_4TLP_STRADDLE(AXISTEN_IF_EXT_512_RC_4TLP_STRADDLE)
   ,.AXISTEN_IF_EXT_512(AXISTEN_IF_EXT_512)
   ,.AXISTEN_IF_CQ_ALIGNMENT_MODE(AXISTEN_IF_CQ_ALIGNMENT_MODE)
   ,.AXISTEN_IF_CC_ALIGNMENT_MODE(AXISTEN_IF_CC_ALIGNMENT_MODE)
   ,.AXISTEN_IF_RQ_ALIGNMENT_MODE(AXISTEN_IF_RQ_ALIGNMENT_MODE)
   ,.AXISTEN_IF_RC_ALIGNMENT_MODE(AXISTEN_IF_RC_ALIGNMENT_MODE)
   ,.AXISTEN_IF_RC_STRADDLE(AXISTEN_IF_RC_STRADDLE)
   ,.AXI4_DATA_WIDTH(AXI4_DATA_WIDTH)
   ,.AXI4_TKEEP_WIDTH(AXI4_TKEEP_WIDTH)
   ,.AXI4_CQ_TUSER_WIDTH(AXI4_CQ_TUSER_WIDTH)
   ,.AXI4_CC_TUSER_WIDTH(AXI4_CC_TUSER_WIDTH)
   ,.AXI4_RQ_TUSER_WIDTH(AXI4_RQ_TUSER_WIDTH)
   ,.AXI4_RC_TUSER_WIDTH(AXI4_RC_TUSER_WIDTH)
   ,.AXI4_CQ_TREADY_WIDTH(AXI4_CQ_TREADY_WIDTH)
   ,.AXI4_CC_TREADY_WIDTH(AXI4_CC_TREADY_WIDTH)
   ,.AXI4_RQ_TREADY_WIDTH(AXI4_RQ_TREADY_WIDTH)
   ,.AXI4_RC_TREADY_WIDTH(AXI4_RC_TREADY_WIDTH)
   ,.AXISTEN_IF_ENABLE_RX_MSG_INTFC(AXISTEN_IF_ENABLE_RX_MSG_INTFC)
   ,.AXISTEN_IF_ENABLE_MSG_ROUTE(AXISTEN_IF_ENABLE_MSG_ROUTE)
   ,.AXISTEN_IF_RX_PARITY_EN(AXISTEN_IF_RX_PARITY_EN)
   ,.AXISTEN_IF_TX_PARITY_EN(AXISTEN_IF_TX_PARITY_EN)
   ,.AXISTEN_IF_ENABLE_CLIENT_TAG(AXISTEN_IF_ENABLE_CLIENT_TAG)
   ,.AXISTEN_IF_ENABLE_256_TAGS(AXISTEN_IF_ENABLE_256_TAGS)
   ,.AXISTEN_IF_COMPL_TIMEOUT_REG0(AXISTEN_IF_COMPL_TIMEOUT_REG0)
   ,.AXISTEN_IF_COMPL_TIMEOUT_REG1(AXISTEN_IF_COMPL_TIMEOUT_REG1)
   ,.AXISTEN_IF_LEGACY_MODE_ENABLE(AXISTEN_IF_LEGACY_MODE_ENABLE)
   ,.AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK(AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK)
   ,.AXISTEN_IF_MSIX_TO_RAM_PIPELINE(AXISTEN_IF_MSIX_TO_RAM_PIPELINE)
   ,.AXISTEN_IF_MSIX_FROM_RAM_PIPELINE(AXISTEN_IF_MSIX_FROM_RAM_PIPELINE)
   ,.AXISTEN_IF_MSIX_RX_PARITY_EN(AXISTEN_IF_MSIX_RX_PARITY_EN)
   ,.AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE(AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE)
   ,.AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT(AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT)
   ,.AXISTEN_IF_CQ_EN_POISONED_MEM_WR(AXISTEN_IF_CQ_EN_POISONED_MEM_WR)
   ,.AXISTEN_IF_RQ_CC_REGISTERED_TREADY(AXISTEN_IF_RQ_CC_REGISTERED_TREADY)
   ,.PM_ASPML0S_TIMEOUT(PM_ASPML0S_TIMEOUT)
   ,.PM_L1_REENTRY_DELAY(PM_L1_REENTRY_DELAY)
   ,.PM_ASPML1_ENTRY_DELAY(PM_ASPML1_ENTRY_DELAY)
   ,.PM_ENABLE_SLOT_POWER_CAPTURE(PM_ENABLE_SLOT_POWER_CAPTURE)
   ,.PM_PME_SERVICE_TIMEOUT_DELAY(PM_PME_SERVICE_TIMEOUT_DELAY)
   ,.PM_PME_TURNOFF_ACK_DELAY(PM_PME_TURNOFF_ACK_DELAY)
   ,.PL_UPSTREAM_FACING(PL_UPSTREAM_FACING)
   ,.PL_LINK_CAP_MAX_LINK_WIDTH(PL_LINK_CAP_MAX_LINK_WIDTH)
   ,.PL_LINK_CAP_MAX_LINK_SPEED(PL_LINK_CAP_MAX_LINK_SPEED)
   ,.PL_DISABLE_DC_BALANCE(PL_DISABLE_DC_BALANCE)
   ,.PL_DISABLE_EI_INFER_IN_L0(PL_DISABLE_EI_INFER_IN_L0)
   ,.PL_N_FTS(PL_N_FTS)
   ,.PL_DISABLE_UPCONFIG_CAPABLE(PL_DISABLE_UPCONFIG_CAPABLE)
   ,.PL_DISABLE_RETRAIN_ON_FRAMING_ERROR(PL_DISABLE_RETRAIN_ON_FRAMING_ERROR)
   ,.PL_DISABLE_RETRAIN_ON_EB_ERROR(PL_DISABLE_RETRAIN_ON_EB_ERROR)
   ,.PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR(PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR)
   ,.PL_REPORT_ALL_PHY_ERRORS(PL_REPORT_ALL_PHY_ERRORS)
   ,.PL_DISABLE_LFSR_UPDATE_ON_SKP(PL_DISABLE_LFSR_UPDATE_ON_SKP)
   ,.PL_LANE0_EQ_CONTROL(PL_LANE0_EQ_CONTROL)
   ,.PL_LANE1_EQ_CONTROL(PL_LANE1_EQ_CONTROL)
   ,.PL_LANE2_EQ_CONTROL(PL_LANE2_EQ_CONTROL)
   ,.PL_LANE3_EQ_CONTROL(PL_LANE3_EQ_CONTROL)
   ,.PL_LANE4_EQ_CONTROL(PL_LANE4_EQ_CONTROL)
   ,.PL_LANE5_EQ_CONTROL(PL_LANE5_EQ_CONTROL)
   ,.PL_LANE6_EQ_CONTROL(PL_LANE6_EQ_CONTROL)
   ,.PL_LANE7_EQ_CONTROL(PL_LANE7_EQ_CONTROL)
   ,.PL_LANE8_EQ_CONTROL(PL_LANE8_EQ_CONTROL)
   ,.PL_LANE9_EQ_CONTROL(PL_LANE9_EQ_CONTROL)
   ,.PL_LANE10_EQ_CONTROL(PL_LANE10_EQ_CONTROL)
   ,.PL_LANE11_EQ_CONTROL(PL_LANE11_EQ_CONTROL)
   ,.PL_LANE12_EQ_CONTROL(PL_LANE12_EQ_CONTROL)
   ,.PL_LANE13_EQ_CONTROL(PL_LANE13_EQ_CONTROL)
   ,.PL_LANE14_EQ_CONTROL(PL_LANE14_EQ_CONTROL)
   ,.PL_LANE15_EQ_CONTROL(PL_LANE15_EQ_CONTROL)
   ,.PL_EQ_BYPASS_PHASE23(PL_EQ_BYPASS_PHASE23)
   ,.PL_EQ_ADAPT_ITER_COUNT(PL_EQ_ADAPT_ITER_COUNT)
   ,.PL_EQ_ADAPT_REJECT_RETRY_COUNT(PL_EQ_ADAPT_REJECT_RETRY_COUNT)
   ,.PL_EQ_SHORT_ADAPT_PHASE(PL_EQ_SHORT_ADAPT_PHASE)
   ,.PL_EQ_ADAPT_DISABLE_COEFF_CHECK(PL_EQ_ADAPT_DISABLE_COEFF_CHECK)
   ,.PL_EQ_ADAPT_DISABLE_PRESET_CHECK(PL_EQ_ADAPT_DISABLE_PRESET_CHECK)
   ,.PL_EQ_DEFAULT_TX_PRESET(PL_EQ_DEFAULT_TX_PRESET)
   ,.PL_EQ_DEFAULT_RX_PRESET_HINT(PL_EQ_DEFAULT_RX_PRESET_HINT)
   ,.PL_EQ_RX_ADAPT_EQ_PHASE0(PL_EQ_RX_ADAPT_EQ_PHASE0)
   ,.PL_EQ_RX_ADAPT_EQ_PHASE1(PL_EQ_RX_ADAPT_EQ_PHASE1)
   ,.PL_EQ_DISABLE_MISMATCH_CHECK(PL_EQ_DISABLE_MISMATCH_CHECK)
   ,.PL_RX_L0S_EXIT_TO_RECOVERY(PL_RX_L0S_EXIT_TO_RECOVERY)
   ,.PL_EQ_TX_8G_EQ_TS2_ENABLE(PL_EQ_TX_8G_EQ_TS2_ENABLE)
   ,.PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4(PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4)
   ,.PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3(PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3)
   ,.PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2(PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2)
   ,.PL_DESKEW_ON_SKIP_IN_GEN12(PL_DESKEW_ON_SKIP_IN_GEN12)
   ,.PL_INFER_EI_DISABLE_REC_RC(PL_INFER_EI_DISABLE_REC_RC)
   ,.PL_INFER_EI_DISABLE_REC_SPD(PL_INFER_EI_DISABLE_REC_SPD)
   ,.PL_INFER_EI_DISABLE_LPBK_ACTIVE(PL_INFER_EI_DISABLE_LPBK_ACTIVE)
   ,.PL_RX_ADAPT_TIMER_RRL_GEN3(PL_RX_ADAPT_TIMER_RRL_GEN3)
   ,.PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS(PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS)
   ,.PL_RX_ADAPT_TIMER_RRL_GEN4(PL_RX_ADAPT_TIMER_RRL_GEN4)
   ,.PL_RX_ADAPT_TIMER_CLWS_GEN3(PL_RX_ADAPT_TIMER_CLWS_GEN3)
   ,.PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS(PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS)
   ,.PL_RX_ADAPT_TIMER_CLWS_GEN4(PL_RX_ADAPT_TIMER_CLWS_GEN4)
   ,.PL_DISABLE_LANE_REVERSAL(PL_DISABLE_LANE_REVERSAL)
   ,.PL_CFG_STATE_ROBUSTNESS_ENABLE(PL_CFG_STATE_ROBUSTNESS_ENABLE)
   ,.PL_REDO_EQ_SOURCE_SELECT(PL_REDO_EQ_SOURCE_SELECT)
   ,.PL_DEEMPH_SOURCE_SELECT(PL_DEEMPH_SOURCE_SELECT)
   ,.PL_EXIT_LOOPBACK_ON_EI_ENTRY(PL_EXIT_LOOPBACK_ON_EI_ENTRY)
   ,.PL_QUIESCE_GUARANTEE_DISABLE(PL_QUIESCE_GUARANTEE_DISABLE)
   ,.PL_SRIS_ENABLE(PL_SRIS_ENABLE)
   ,.PL_SRIS_SKPOS_GEN_SPD_VEC(PL_SRIS_SKPOS_GEN_SPD_VEC)
   ,.PL_SRIS_SKPOS_REC_SPD_VEC(PL_SRIS_SKPOS_REC_SPD_VEC)
   ,.PL_SIM_FAST_LINK_TRAINING(PL_SIM_FAST_LINK_TRAINING)
   ,.PL_USER_SPARE(PL_USER_SPARE)
   ,.LL_ACK_TIMEOUT_EN(LL_ACK_TIMEOUT_EN)
   ,.LL_ACK_TIMEOUT(LL_ACK_TIMEOUT)
   ,.LL_ACK_TIMEOUT_FUNC(LL_ACK_TIMEOUT_FUNC)
   ,.LL_REPLAY_TIMEOUT_EN(LL_REPLAY_TIMEOUT_EN)
   ,.LL_REPLAY_TIMEOUT(LL_REPLAY_TIMEOUT)
   ,.LL_REPLAY_TIMEOUT_FUNC(LL_REPLAY_TIMEOUT_FUNC)
   ,.LL_REPLAY_TO_RAM_PIPELINE(LL_REPLAY_TO_RAM_PIPELINE)
   ,.LL_REPLAY_FROM_RAM_PIPELINE(LL_REPLAY_FROM_RAM_PIPELINE)
   ,.LL_DISABLE_SCHED_TX_NAK(LL_DISABLE_SCHED_TX_NAK)
   ,.LL_TX_TLP_PARITY_CHK(LL_TX_TLP_PARITY_CHK)
   ,.LL_RX_TLP_PARITY_GEN(LL_RX_TLP_PARITY_GEN)
   ,.LL_USER_SPARE(LL_USER_SPARE)
   ,.IS_SWITCH_PORT(IS_SWITCH_PORT)
   ,.CFG_BYPASS_MODE_ENABLE(CFG_BYPASS_MODE_ENABLE)
   ,.TL_PF_ENABLE_REG(TL_PF_ENABLE_REG)
   ,.TL_CREDITS_CD(TL_CREDITS_CD)
   ,.TL_CREDITS_CH(TL_CREDITS_CH)
   ,.TL_COMPLETION_RAM_SIZE(TL_COMPLETION_RAM_SIZE)
   ,.TL_COMPLETION_RAM_NUM_TLPS(TL_COMPLETION_RAM_NUM_TLPS)
   ,.TL_CREDITS_NPD(TL_CREDITS_NPD)
   ,.TL_CREDITS_NPH(TL_CREDITS_NPH)
   ,.TL_CREDITS_PD(TL_CREDITS_PD)
   ,.TL_CREDITS_PH(TL_CREDITS_PH)
   ,.TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE(TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE)
   ,.TL_RX_COMPLETION_TO_RAM_READ_PIPELINE(TL_RX_COMPLETION_TO_RAM_READ_PIPELINE)
   ,.TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE(TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE)
   ,.TL_POSTED_RAM_SIZE(TL_POSTED_RAM_SIZE)
   ,.TL_RX_POSTED_TO_RAM_WRITE_PIPELINE(TL_RX_POSTED_TO_RAM_WRITE_PIPELINE)
   ,.TL_RX_POSTED_TO_RAM_READ_PIPELINE(TL_RX_POSTED_TO_RAM_READ_PIPELINE)
   ,.TL_RX_POSTED_FROM_RAM_READ_PIPELINE(TL_RX_POSTED_FROM_RAM_READ_PIPELINE)
   ,.TL_TX_MUX_STRICT_PRIORITY(TL_TX_MUX_STRICT_PRIORITY)
   ,.TL_TX_TLP_STRADDLE_ENABLE(TL_TX_TLP_STRADDLE_ENABLE)
   ,.TL_TX_TLP_TERMINATE_PARITY(TL_TX_TLP_TERMINATE_PARITY)
   ,.TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT(TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT)
   ,.TL_FC_UPDATE_MIN_INTERVAL_TIME(TL_FC_UPDATE_MIN_INTERVAL_TIME)
   ,.TL_USER_SPARE(TL_USER_SPARE)
   ,.PF0_CLASS_CODE(PF0_CLASS_CODE)
   ,.PF1_CLASS_CODE(PF1_CLASS_CODE)
   ,.PF2_CLASS_CODE(PF2_CLASS_CODE)
   ,.PF3_CLASS_CODE(PF3_CLASS_CODE)
   ,.PF0_INTERRUPT_PIN(PF0_INTERRUPT_PIN)
   ,.PF1_INTERRUPT_PIN(PF1_INTERRUPT_PIN)
   ,.PF2_INTERRUPT_PIN(PF2_INTERRUPT_PIN)
   ,.PF3_INTERRUPT_PIN(PF3_INTERRUPT_PIN)
   ,.PF0_CAPABILITY_POINTER(PF0_CAPABILITY_POINTER)
   ,.PF1_CAPABILITY_POINTER(PF1_CAPABILITY_POINTER)
   ,.PF2_CAPABILITY_POINTER(PF2_CAPABILITY_POINTER)
   ,.PF3_CAPABILITY_POINTER(PF3_CAPABILITY_POINTER)
   ,.VF0_CAPABILITY_POINTER(VF0_CAPABILITY_POINTER)
   ,.LEGACY_CFG_EXTEND_INTERFACE_ENABLE(LEGACY_CFG_EXTEND_INTERFACE_ENABLE)
   ,.EXTENDED_CFG_EXTEND_INTERFACE_ENABLE(EXTENDED_CFG_EXTEND_INTERFACE_ENABLE)
   ,.TL2CFG_IF_PARITY_CHK(TL2CFG_IF_PARITY_CHK)
   ,.HEADER_TYPE_OVERRIDE(HEADER_TYPE_OVERRIDE)
   ,.PF0_BAR0_CONTROL(PF0_BAR0_CONTROL)
   ,.PF1_BAR0_CONTROL(PF1_BAR0_CONTROL)
   ,.PF2_BAR0_CONTROL(PF2_BAR0_CONTROL)
   ,.PF3_BAR0_CONTROL(PF3_BAR0_CONTROL)
   ,.PF0_BAR0_APERTURE_SIZE(PF0_BAR0_APERTURE_SIZE)
   ,.PF1_BAR0_APERTURE_SIZE(PF1_BAR0_APERTURE_SIZE)
   ,.PF2_BAR0_APERTURE_SIZE(PF2_BAR0_APERTURE_SIZE)
   ,.PF3_BAR0_APERTURE_SIZE(PF3_BAR0_APERTURE_SIZE)
   ,.PF0_BAR1_CONTROL(PF0_BAR1_CONTROL)
   ,.PF1_BAR1_CONTROL(PF1_BAR1_CONTROL)
   ,.PF2_BAR1_CONTROL(PF2_BAR1_CONTROL)
   ,.PF3_BAR1_CONTROL(PF3_BAR1_CONTROL)
   ,.PF0_BAR1_APERTURE_SIZE(PF0_BAR1_APERTURE_SIZE)
   ,.PF1_BAR1_APERTURE_SIZE(PF1_BAR1_APERTURE_SIZE)
   ,.PF2_BAR1_APERTURE_SIZE(PF2_BAR1_APERTURE_SIZE)
   ,.PF3_BAR1_APERTURE_SIZE(PF3_BAR1_APERTURE_SIZE)
   ,.PF0_BAR2_CONTROL(PF0_BAR2_CONTROL)
   ,.PF1_BAR2_CONTROL(PF1_BAR2_CONTROL)
   ,.PF2_BAR2_CONTROL(PF2_BAR2_CONTROL)
   ,.PF3_BAR2_CONTROL(PF3_BAR2_CONTROL)
   ,.PF0_BAR2_APERTURE_SIZE(PF0_BAR2_APERTURE_SIZE)
   ,.PF1_BAR2_APERTURE_SIZE(PF1_BAR2_APERTURE_SIZE)
   ,.PF2_BAR2_APERTURE_SIZE(PF2_BAR2_APERTURE_SIZE)
   ,.PF3_BAR2_APERTURE_SIZE(PF3_BAR2_APERTURE_SIZE)
   ,.PF0_BAR3_CONTROL(PF0_BAR3_CONTROL)
   ,.PF1_BAR3_CONTROL(PF1_BAR3_CONTROL)
   ,.PF2_BAR3_CONTROL(PF2_BAR3_CONTROL)
   ,.PF3_BAR3_CONTROL(PF3_BAR3_CONTROL)
   ,.PF0_BAR3_APERTURE_SIZE(PF0_BAR3_APERTURE_SIZE)
   ,.PF1_BAR3_APERTURE_SIZE(PF1_BAR3_APERTURE_SIZE)
   ,.PF2_BAR3_APERTURE_SIZE(PF2_BAR3_APERTURE_SIZE)
   ,.PF3_BAR3_APERTURE_SIZE(PF3_BAR3_APERTURE_SIZE)
   ,.PF0_BAR4_CONTROL(PF0_BAR4_CONTROL)
   ,.PF1_BAR4_CONTROL(PF1_BAR4_CONTROL)
   ,.PF2_BAR4_CONTROL(PF2_BAR4_CONTROL)
   ,.PF3_BAR4_CONTROL(PF3_BAR4_CONTROL)
   ,.PF0_BAR4_APERTURE_SIZE(PF0_BAR4_APERTURE_SIZE)
   ,.PF1_BAR4_APERTURE_SIZE(PF1_BAR4_APERTURE_SIZE)
   ,.PF2_BAR4_APERTURE_SIZE(PF2_BAR4_APERTURE_SIZE)
   ,.PF3_BAR4_APERTURE_SIZE(PF3_BAR4_APERTURE_SIZE)
   ,.PF0_BAR5_CONTROL(PF0_BAR5_CONTROL)
   ,.PF1_BAR5_CONTROL(PF1_BAR5_CONTROL)
   ,.PF2_BAR5_CONTROL(PF2_BAR5_CONTROL)
   ,.PF3_BAR5_CONTROL(PF3_BAR5_CONTROL)
   ,.PF0_BAR5_APERTURE_SIZE(PF0_BAR5_APERTURE_SIZE)
   ,.PF1_BAR5_APERTURE_SIZE(PF1_BAR5_APERTURE_SIZE)
   ,.PF2_BAR5_APERTURE_SIZE(PF2_BAR5_APERTURE_SIZE)
   ,.PF3_BAR5_APERTURE_SIZE(PF3_BAR5_APERTURE_SIZE)
   ,.PF0_EXPANSION_ROM_ENABLE(PF0_EXPANSION_ROM_ENABLE)
   ,.PF1_EXPANSION_ROM_ENABLE(PF1_EXPANSION_ROM_ENABLE)
   ,.PF2_EXPANSION_ROM_ENABLE(PF2_EXPANSION_ROM_ENABLE)
   ,.PF3_EXPANSION_ROM_ENABLE(PF3_EXPANSION_ROM_ENABLE)
   ,.PF0_EXPANSION_ROM_APERTURE_SIZE(PF0_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF1_EXPANSION_ROM_APERTURE_SIZE(PF1_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF2_EXPANSION_ROM_APERTURE_SIZE(PF2_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF3_EXPANSION_ROM_APERTURE_SIZE(PF3_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF0_PCIE_CAP_NEXTPTR(PF0_PCIE_CAP_NEXTPTR)
   ,.PF1_PCIE_CAP_NEXTPTR(PF1_PCIE_CAP_NEXTPTR)
   ,.PF2_PCIE_CAP_NEXTPTR(PF2_PCIE_CAP_NEXTPTR)
   ,.PF3_PCIE_CAP_NEXTPTR(PF3_PCIE_CAP_NEXTPTR)
   ,.VFG0_PCIE_CAP_NEXTPTR(VFG0_PCIE_CAP_NEXTPTR)
   ,.VFG1_PCIE_CAP_NEXTPTR(VFG1_PCIE_CAP_NEXTPTR)
   ,.VFG2_PCIE_CAP_NEXTPTR(VFG2_PCIE_CAP_NEXTPTR)
   ,.VFG3_PCIE_CAP_NEXTPTR(VFG3_PCIE_CAP_NEXTPTR)
   ,.PF0_DEV_CAP_MAX_PAYLOAD_SIZE(PF0_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF1_DEV_CAP_MAX_PAYLOAD_SIZE(PF1_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF2_DEV_CAP_MAX_PAYLOAD_SIZE(PF2_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF3_DEV_CAP_MAX_PAYLOAD_SIZE(PF3_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF0_DEV_CAP_EXT_TAG_SUPPORTED(PF0_DEV_CAP_EXT_TAG_SUPPORTED)
   ,.PF0_DEV_CAP_ENDPOINT_L0S_LATENCY(PF0_DEV_CAP_ENDPOINT_L0S_LATENCY)
   ,.PF0_DEV_CAP_ENDPOINT_L1_LATENCY(PF0_DEV_CAP_ENDPOINT_L1_LATENCY)
   ,.PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE(PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE)
   ,.PF0_LINK_CAP_ASPM_SUPPORT(PF0_LINK_CAP_ASPM_SUPPORT)
   ,.PF0_LINK_CONTROL_RCB(PF0_LINK_CONTROL_RCB)
   ,.PF0_LINK_STATUS_SLOT_CLOCK_CONFIG(PF0_LINK_STATUS_SLOT_CLOCK_CONFIG)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4)
   ,.PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE(PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE)
   ,.PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT(PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT(PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT(PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_LTR_SUPPORT(PF0_DEV_CAP2_LTR_SUPPORT)
   ,.PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT(PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_OBFF_SUPPORT(PF0_DEV_CAP2_OBFF_SUPPORT)
   ,.PF0_DEV_CAP2_ARI_FORWARD_ENABLE(PF0_DEV_CAP2_ARI_FORWARD_ENABLE)
   ,.PF0_MSI_CAP_NEXTPTR(PF0_MSI_CAP_NEXTPTR)
   ,.PF1_MSI_CAP_NEXTPTR(PF1_MSI_CAP_NEXTPTR)
   ,.PF2_MSI_CAP_NEXTPTR(PF2_MSI_CAP_NEXTPTR)
   ,.PF3_MSI_CAP_NEXTPTR(PF3_MSI_CAP_NEXTPTR)
   ,.PF0_MSI_CAP_PERVECMASKCAP(PF0_MSI_CAP_PERVECMASKCAP)
   ,.PF1_MSI_CAP_PERVECMASKCAP(PF1_MSI_CAP_PERVECMASKCAP)
   ,.PF2_MSI_CAP_PERVECMASKCAP(PF2_MSI_CAP_PERVECMASKCAP)
   ,.PF3_MSI_CAP_PERVECMASKCAP(PF3_MSI_CAP_PERVECMASKCAP)
   ,.PF0_MSI_CAP_MULTIMSGCAP(PF0_MSI_CAP_MULTIMSGCAP)
   ,.PF1_MSI_CAP_MULTIMSGCAP(PF1_MSI_CAP_MULTIMSGCAP)
   ,.PF2_MSI_CAP_MULTIMSGCAP(PF2_MSI_CAP_MULTIMSGCAP)
   ,.PF3_MSI_CAP_MULTIMSGCAP(PF3_MSI_CAP_MULTIMSGCAP)
   ,.PF0_MSIX_CAP_NEXTPTR(PF0_MSIX_CAP_NEXTPTR)
   ,.PF1_MSIX_CAP_NEXTPTR(PF1_MSIX_CAP_NEXTPTR)
   ,.PF2_MSIX_CAP_NEXTPTR(PF2_MSIX_CAP_NEXTPTR)
   ,.PF3_MSIX_CAP_NEXTPTR(PF3_MSIX_CAP_NEXTPTR)
   ,.VFG0_MSIX_CAP_NEXTPTR(VFG0_MSIX_CAP_NEXTPTR)
   ,.VFG1_MSIX_CAP_NEXTPTR(VFG1_MSIX_CAP_NEXTPTR)
   ,.VFG2_MSIX_CAP_NEXTPTR(VFG2_MSIX_CAP_NEXTPTR)
   ,.VFG3_MSIX_CAP_NEXTPTR(VFG3_MSIX_CAP_NEXTPTR)
   ,.PF0_MSIX_CAP_PBA_BIR(PF0_MSIX_CAP_PBA_BIR)
   ,.PF1_MSIX_CAP_PBA_BIR(PF1_MSIX_CAP_PBA_BIR)
   ,.PF2_MSIX_CAP_PBA_BIR(PF2_MSIX_CAP_PBA_BIR)
   ,.PF3_MSIX_CAP_PBA_BIR(PF3_MSIX_CAP_PBA_BIR)
   ,.VFG0_MSIX_CAP_PBA_BIR(VFG0_MSIX_CAP_PBA_BIR)
   ,.VFG1_MSIX_CAP_PBA_BIR(VFG1_MSIX_CAP_PBA_BIR)
   ,.VFG2_MSIX_CAP_PBA_BIR(VFG2_MSIX_CAP_PBA_BIR)
   ,.VFG3_MSIX_CAP_PBA_BIR(VFG3_MSIX_CAP_PBA_BIR)
   ,.PF0_MSIX_CAP_PBA_OFFSET(PF0_MSIX_CAP_PBA_OFFSET)
   ,.PF1_MSIX_CAP_PBA_OFFSET(PF1_MSIX_CAP_PBA_OFFSET)
   ,.PF2_MSIX_CAP_PBA_OFFSET(PF2_MSIX_CAP_PBA_OFFSET)
   ,.PF3_MSIX_CAP_PBA_OFFSET(PF3_MSIX_CAP_PBA_OFFSET)
   ,.VFG0_MSIX_CAP_PBA_OFFSET(VFG0_MSIX_CAP_PBA_OFFSET)
   ,.VFG1_MSIX_CAP_PBA_OFFSET(VFG1_MSIX_CAP_PBA_OFFSET)
   ,.VFG2_MSIX_CAP_PBA_OFFSET(VFG2_MSIX_CAP_PBA_OFFSET)
   ,.VFG3_MSIX_CAP_PBA_OFFSET(VFG3_MSIX_CAP_PBA_OFFSET)
   ,.PF0_MSIX_CAP_TABLE_BIR(PF0_MSIX_CAP_TABLE_BIR)
   ,.PF1_MSIX_CAP_TABLE_BIR(PF1_MSIX_CAP_TABLE_BIR)
   ,.PF2_MSIX_CAP_TABLE_BIR(PF2_MSIX_CAP_TABLE_BIR)
   ,.PF3_MSIX_CAP_TABLE_BIR(PF3_MSIX_CAP_TABLE_BIR)
   ,.VFG0_MSIX_CAP_TABLE_BIR(VFG0_MSIX_CAP_TABLE_BIR)
   ,.VFG1_MSIX_CAP_TABLE_BIR(VFG1_MSIX_CAP_TABLE_BIR)
   ,.VFG2_MSIX_CAP_TABLE_BIR(VFG2_MSIX_CAP_TABLE_BIR)
   ,.VFG3_MSIX_CAP_TABLE_BIR(VFG3_MSIX_CAP_TABLE_BIR)
   ,.PF0_MSIX_CAP_TABLE_OFFSET(PF0_MSIX_CAP_TABLE_OFFSET)
   ,.PF1_MSIX_CAP_TABLE_OFFSET(PF1_MSIX_CAP_TABLE_OFFSET)
   ,.PF2_MSIX_CAP_TABLE_OFFSET(PF2_MSIX_CAP_TABLE_OFFSET)
   ,.PF3_MSIX_CAP_TABLE_OFFSET(PF3_MSIX_CAP_TABLE_OFFSET)
   ,.VFG0_MSIX_CAP_TABLE_OFFSET(VFG0_MSIX_CAP_TABLE_OFFSET)
   ,.VFG1_MSIX_CAP_TABLE_OFFSET(VFG1_MSIX_CAP_TABLE_OFFSET)
   ,.VFG2_MSIX_CAP_TABLE_OFFSET(VFG2_MSIX_CAP_TABLE_OFFSET)
   ,.VFG3_MSIX_CAP_TABLE_OFFSET(VFG3_MSIX_CAP_TABLE_OFFSET)
   ,.PF0_MSIX_CAP_TABLE_SIZE(PF0_MSIX_CAP_TABLE_SIZE)
   ,.PF1_MSIX_CAP_TABLE_SIZE(PF1_MSIX_CAP_TABLE_SIZE)
   ,.PF2_MSIX_CAP_TABLE_SIZE(PF2_MSIX_CAP_TABLE_SIZE)
   ,.PF3_MSIX_CAP_TABLE_SIZE(PF3_MSIX_CAP_TABLE_SIZE)
   ,.VFG0_MSIX_CAP_TABLE_SIZE(VFG0_MSIX_CAP_TABLE_SIZE)
   ,.VFG1_MSIX_CAP_TABLE_SIZE(VFG1_MSIX_CAP_TABLE_SIZE)
   ,.VFG2_MSIX_CAP_TABLE_SIZE(VFG2_MSIX_CAP_TABLE_SIZE)
   ,.VFG3_MSIX_CAP_TABLE_SIZE(VFG3_MSIX_CAP_TABLE_SIZE)
   ,.PF0_MSIX_VECTOR_COUNT(PF0_MSIX_VECTOR_COUNT)
   ,.PF0_PM_CAP_ID(PF0_PM_CAP_ID)
   ,.PF0_PM_CAP_NEXTPTR(PF0_PM_CAP_NEXTPTR)
   ,.PF1_PM_CAP_NEXTPTR(PF1_PM_CAP_NEXTPTR)
   ,.PF2_PM_CAP_NEXTPTR(PF2_PM_CAP_NEXTPTR)
   ,.PF3_PM_CAP_NEXTPTR(PF3_PM_CAP_NEXTPTR)
   ,.PF0_PM_CAP_PMESUPPORT_D3HOT(PF0_PM_CAP_PMESUPPORT_D3HOT)
   ,.PF0_PM_CAP_PMESUPPORT_D1(PF0_PM_CAP_PMESUPPORT_D1)
   ,.PF0_PM_CAP_PMESUPPORT_D0(PF0_PM_CAP_PMESUPPORT_D0)
   ,.PF0_PM_CAP_SUPP_D1_STATE(PF0_PM_CAP_SUPP_D1_STATE)
   ,.PF0_PM_CAP_VER_ID(PF0_PM_CAP_VER_ID)
   ,.PF0_PM_CSR_NOSOFTRESET(PF0_PM_CSR_NOSOFTRESET)
   ,.PM_ENABLE_L23_ENTRY(PM_ENABLE_L23_ENTRY)
   ,.DNSTREAM_LINK_NUM(DNSTREAM_LINK_NUM)
   ,.AUTO_FLR_RESPONSE(AUTO_FLR_RESPONSE)
   ,.PF0_DSN_CAP_NEXTPTR(PF0_DSN_CAP_NEXTPTR)
   ,.PF1_DSN_CAP_NEXTPTR(PF1_DSN_CAP_NEXTPTR)
   ,.PF2_DSN_CAP_NEXTPTR(PF2_DSN_CAP_NEXTPTR)
   ,.PF3_DSN_CAP_NEXTPTR(PF3_DSN_CAP_NEXTPTR)
   ,.DSN_CAP_ENABLE(DSN_CAP_ENABLE)
   ,.PF0_VC_CAP_VER(PF0_VC_CAP_VER)
   ,.PF0_VC_CAP_NEXTPTR(PF0_VC_CAP_NEXTPTR)
   ,.PF0_VC_CAP_ENABLE(PF0_VC_CAP_ENABLE)
   ,.PF0_SECONDARY_PCIE_CAP_NEXTPTR(PF0_SECONDARY_PCIE_CAP_NEXTPTR)
   ,.PF0_AER_CAP_NEXTPTR(PF0_AER_CAP_NEXTPTR)
   ,.PF1_AER_CAP_NEXTPTR(PF1_AER_CAP_NEXTPTR)
   ,.PF2_AER_CAP_NEXTPTR(PF2_AER_CAP_NEXTPTR)
   ,.PF3_AER_CAP_NEXTPTR(PF3_AER_CAP_NEXTPTR)
   ,.PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE(PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE)
   ,.ARI_CAP_ENABLE(ARI_CAP_ENABLE)
   ,.PF0_ARI_CAP_NEXTPTR(PF0_ARI_CAP_NEXTPTR)
   ,.PF1_ARI_CAP_NEXTPTR(PF1_ARI_CAP_NEXTPTR)
   ,.PF2_ARI_CAP_NEXTPTR(PF2_ARI_CAP_NEXTPTR)
   ,.PF3_ARI_CAP_NEXTPTR(PF3_ARI_CAP_NEXTPTR)
   ,.VFG0_ARI_CAP_NEXTPTR(VFG0_ARI_CAP_NEXTPTR)
   ,.VFG1_ARI_CAP_NEXTPTR(VFG1_ARI_CAP_NEXTPTR)
   ,.VFG2_ARI_CAP_NEXTPTR(VFG2_ARI_CAP_NEXTPTR)
   ,.VFG3_ARI_CAP_NEXTPTR(VFG3_ARI_CAP_NEXTPTR)
   ,.PF0_ARI_CAP_VER(PF0_ARI_CAP_VER)
   ,.PF0_ARI_CAP_NEXT_FUNC(PF0_ARI_CAP_NEXT_FUNC)
   ,.PF1_ARI_CAP_NEXT_FUNC(PF1_ARI_CAP_NEXT_FUNC)
   ,.PF2_ARI_CAP_NEXT_FUNC(PF2_ARI_CAP_NEXT_FUNC)
   ,.PF3_ARI_CAP_NEXT_FUNC(PF3_ARI_CAP_NEXT_FUNC)
   ,.PF0_LTR_CAP_NEXTPTR(PF0_LTR_CAP_NEXTPTR)
   ,.PF0_LTR_CAP_VER(PF0_LTR_CAP_VER)
   ,.PF0_LTR_CAP_MAX_SNOOP_LAT(PF0_LTR_CAP_MAX_SNOOP_LAT)
   ,.PF0_LTR_CAP_MAX_NOSNOOP_LAT(PF0_LTR_CAP_MAX_NOSNOOP_LAT)
   ,.LTR_TX_MESSAGE_ON_LTR_ENABLE(LTR_TX_MESSAGE_ON_LTR_ENABLE)
   ,.LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE(LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE)
   ,.LTR_TX_MESSAGE_MINIMUM_INTERVAL(LTR_TX_MESSAGE_MINIMUM_INTERVAL)
   ,.SRIOV_CAP_ENABLE(SRIOV_CAP_ENABLE)
   ,.PF0_SRIOV_CAP_NEXTPTR(PF0_SRIOV_CAP_NEXTPTR)
   ,.PF1_SRIOV_CAP_NEXTPTR(PF1_SRIOV_CAP_NEXTPTR)
   ,.PF2_SRIOV_CAP_NEXTPTR(PF2_SRIOV_CAP_NEXTPTR)
   ,.PF3_SRIOV_CAP_NEXTPTR(PF3_SRIOV_CAP_NEXTPTR)
   ,.PF0_SRIOV_CAP_VER(PF0_SRIOV_CAP_VER)
   ,.PF1_SRIOV_CAP_VER(PF1_SRIOV_CAP_VER)
   ,.PF2_SRIOV_CAP_VER(PF2_SRIOV_CAP_VER)
   ,.PF3_SRIOV_CAP_VER(PF3_SRIOV_CAP_VER)
   ,.PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF0_SRIOV_CAP_INITIAL_VF(PF0_SRIOV_CAP_INITIAL_VF)
   ,.PF1_SRIOV_CAP_INITIAL_VF(PF1_SRIOV_CAP_INITIAL_VF)
   ,.PF2_SRIOV_CAP_INITIAL_VF(PF2_SRIOV_CAP_INITIAL_VF)
   ,.PF3_SRIOV_CAP_INITIAL_VF(PF3_SRIOV_CAP_INITIAL_VF)
   ,.PF0_SRIOV_CAP_TOTAL_VF(PF0_SRIOV_CAP_TOTAL_VF)
   ,.PF1_SRIOV_CAP_TOTAL_VF(PF1_SRIOV_CAP_TOTAL_VF)
   ,.PF2_SRIOV_CAP_TOTAL_VF(PF2_SRIOV_CAP_TOTAL_VF)
   ,.PF3_SRIOV_CAP_TOTAL_VF(PF3_SRIOV_CAP_TOTAL_VF)
   ,.PF0_SRIOV_FUNC_DEP_LINK(PF0_SRIOV_FUNC_DEP_LINK)
   ,.PF1_SRIOV_FUNC_DEP_LINK(PF1_SRIOV_FUNC_DEP_LINK)
   ,.PF2_SRIOV_FUNC_DEP_LINK(PF2_SRIOV_FUNC_DEP_LINK)
   ,.PF3_SRIOV_FUNC_DEP_LINK(PF3_SRIOV_FUNC_DEP_LINK)
   ,.PF0_SRIOV_FIRST_VF_OFFSET(PF0_SRIOV_FIRST_VF_OFFSET)
   ,.PF1_SRIOV_FIRST_VF_OFFSET(PF1_SRIOV_FIRST_VF_OFFSET)
   ,.PF2_SRIOV_FIRST_VF_OFFSET(PF2_SRIOV_FIRST_VF_OFFSET)
   ,.PF3_SRIOV_FIRST_VF_OFFSET(PF3_SRIOV_FIRST_VF_OFFSET)
   ,.PF0_SRIOV_VF_DEVICE_ID(PF0_SRIOV_VF_DEVICE_ID)
   ,.PF1_SRIOV_VF_DEVICE_ID(PF1_SRIOV_VF_DEVICE_ID)
   ,.PF2_SRIOV_VF_DEVICE_ID(PF2_SRIOV_VF_DEVICE_ID)
   ,.PF3_SRIOV_VF_DEVICE_ID(PF3_SRIOV_VF_DEVICE_ID)
   ,.PF0_SRIOV_SUPPORTED_PAGE_SIZE(PF0_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF1_SRIOV_SUPPORTED_PAGE_SIZE(PF1_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF2_SRIOV_SUPPORTED_PAGE_SIZE(PF2_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF3_SRIOV_SUPPORTED_PAGE_SIZE(PF3_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF0_SRIOV_BAR0_CONTROL(PF0_SRIOV_BAR0_CONTROL)
   ,.PF1_SRIOV_BAR0_CONTROL(PF1_SRIOV_BAR0_CONTROL)
   ,.PF2_SRIOV_BAR0_CONTROL(PF2_SRIOV_BAR0_CONTROL)
   ,.PF3_SRIOV_BAR0_CONTROL(PF3_SRIOV_BAR0_CONTROL)
   ,.PF0_SRIOV_BAR0_APERTURE_SIZE(PF0_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR0_APERTURE_SIZE(PF1_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR0_APERTURE_SIZE(PF2_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR0_APERTURE_SIZE(PF3_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR1_CONTROL(PF0_SRIOV_BAR1_CONTROL)
   ,.PF1_SRIOV_BAR1_CONTROL(PF1_SRIOV_BAR1_CONTROL)
   ,.PF2_SRIOV_BAR1_CONTROL(PF2_SRIOV_BAR1_CONTROL)
   ,.PF3_SRIOV_BAR1_CONTROL(PF3_SRIOV_BAR1_CONTROL)
   ,.PF0_SRIOV_BAR1_APERTURE_SIZE(PF0_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR1_APERTURE_SIZE(PF1_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR1_APERTURE_SIZE(PF2_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR1_APERTURE_SIZE(PF3_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR2_CONTROL(PF0_SRIOV_BAR2_CONTROL)
   ,.PF1_SRIOV_BAR2_CONTROL(PF1_SRIOV_BAR2_CONTROL)
   ,.PF2_SRIOV_BAR2_CONTROL(PF2_SRIOV_BAR2_CONTROL)
   ,.PF3_SRIOV_BAR2_CONTROL(PF3_SRIOV_BAR2_CONTROL)
   ,.PF0_SRIOV_BAR2_APERTURE_SIZE(PF0_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR2_APERTURE_SIZE(PF1_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR2_APERTURE_SIZE(PF2_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR2_APERTURE_SIZE(PF3_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR3_CONTROL(PF0_SRIOV_BAR3_CONTROL)
   ,.PF1_SRIOV_BAR3_CONTROL(PF1_SRIOV_BAR3_CONTROL)
   ,.PF2_SRIOV_BAR3_CONTROL(PF2_SRIOV_BAR3_CONTROL)
   ,.PF3_SRIOV_BAR3_CONTROL(PF3_SRIOV_BAR3_CONTROL)
   ,.PF0_SRIOV_BAR3_APERTURE_SIZE(PF0_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR3_APERTURE_SIZE(PF1_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR3_APERTURE_SIZE(PF2_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR3_APERTURE_SIZE(PF3_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR4_CONTROL(PF0_SRIOV_BAR4_CONTROL)
   ,.PF1_SRIOV_BAR4_CONTROL(PF1_SRIOV_BAR4_CONTROL)
   ,.PF2_SRIOV_BAR4_CONTROL(PF2_SRIOV_BAR4_CONTROL)
   ,.PF3_SRIOV_BAR4_CONTROL(PF3_SRIOV_BAR4_CONTROL)
   ,.PF0_SRIOV_BAR4_APERTURE_SIZE(PF0_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR4_APERTURE_SIZE(PF1_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR4_APERTURE_SIZE(PF2_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR4_APERTURE_SIZE(PF3_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR5_CONTROL(PF0_SRIOV_BAR5_CONTROL)
   ,.PF1_SRIOV_BAR5_CONTROL(PF1_SRIOV_BAR5_CONTROL)
   ,.PF2_SRIOV_BAR5_CONTROL(PF2_SRIOV_BAR5_CONTROL)
   ,.PF3_SRIOV_BAR5_CONTROL(PF3_SRIOV_BAR5_CONTROL)
   ,.PF0_SRIOV_BAR5_APERTURE_SIZE(PF0_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR5_APERTURE_SIZE(PF1_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR5_APERTURE_SIZE(PF2_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR5_APERTURE_SIZE(PF3_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF0_TPHR_CAP_NEXTPTR(PF0_TPHR_CAP_NEXTPTR)
   ,.PF1_TPHR_CAP_NEXTPTR(PF1_TPHR_CAP_NEXTPTR)
   ,.PF2_TPHR_CAP_NEXTPTR(PF2_TPHR_CAP_NEXTPTR)
   ,.PF3_TPHR_CAP_NEXTPTR(PF3_TPHR_CAP_NEXTPTR)
   ,.VFG0_TPHR_CAP_NEXTPTR(VFG0_TPHR_CAP_NEXTPTR)
   ,.VFG1_TPHR_CAP_NEXTPTR(VFG1_TPHR_CAP_NEXTPTR)
   ,.VFG2_TPHR_CAP_NEXTPTR(VFG2_TPHR_CAP_NEXTPTR)
   ,.VFG3_TPHR_CAP_NEXTPTR(VFG3_TPHR_CAP_NEXTPTR)
   ,.PF0_TPHR_CAP_VER(PF0_TPHR_CAP_VER)
   ,.PF0_TPHR_CAP_INT_VEC_MODE(PF0_TPHR_CAP_INT_VEC_MODE)
   ,.PF0_TPHR_CAP_DEV_SPECIFIC_MODE(PF0_TPHR_CAP_DEV_SPECIFIC_MODE)
   ,.PF0_TPHR_CAP_ST_TABLE_LOC(PF0_TPHR_CAP_ST_TABLE_LOC)
   ,.PF0_TPHR_CAP_ST_TABLE_SIZE(PF0_TPHR_CAP_ST_TABLE_SIZE)
   ,.PF0_TPHR_CAP_ST_MODE_SEL(PF0_TPHR_CAP_ST_MODE_SEL)
   ,.PF1_TPHR_CAP_ST_MODE_SEL(PF1_TPHR_CAP_ST_MODE_SEL)
   ,.PF2_TPHR_CAP_ST_MODE_SEL(PF2_TPHR_CAP_ST_MODE_SEL)
   ,.PF3_TPHR_CAP_ST_MODE_SEL(PF3_TPHR_CAP_ST_MODE_SEL)
   ,.VFG0_TPHR_CAP_ST_MODE_SEL(VFG0_TPHR_CAP_ST_MODE_SEL)
   ,.VFG1_TPHR_CAP_ST_MODE_SEL(VFG1_TPHR_CAP_ST_MODE_SEL)
   ,.VFG2_TPHR_CAP_ST_MODE_SEL(VFG2_TPHR_CAP_ST_MODE_SEL)
   ,.VFG3_TPHR_CAP_ST_MODE_SEL(VFG3_TPHR_CAP_ST_MODE_SEL)
   ,.PF0_TPHR_CAP_ENABLE(PF0_TPHR_CAP_ENABLE)
   ,.TPH_TO_RAM_PIPELINE(TPH_TO_RAM_PIPELINE)
   ,.TPH_FROM_RAM_PIPELINE(TPH_FROM_RAM_PIPELINE)
   ,.MCAP_ENABLE(MCAP_ENABLE)
   ,.MCAP_CONFIGURE_OVERRIDE(MCAP_CONFIGURE_OVERRIDE)
   ,.MCAP_CAP_NEXTPTR(MCAP_CAP_NEXTPTR)
   ,.MCAP_VSEC_ID(MCAP_VSEC_ID)
   ,.MCAP_VSEC_REV(MCAP_VSEC_REV)
   ,.MCAP_VSEC_LEN(MCAP_VSEC_LEN)
   ,.MCAP_FPGA_BITSTREAM_VERSION(MCAP_FPGA_BITSTREAM_VERSION)
   ,.MCAP_INTERRUPT_ON_MCAP_EOS(MCAP_INTERRUPT_ON_MCAP_EOS)
   ,.MCAP_INTERRUPT_ON_MCAP_ERROR(MCAP_INTERRUPT_ON_MCAP_ERROR)
   ,.MCAP_INPUT_GATE_DESIGN_SWITCH(MCAP_INPUT_GATE_DESIGN_SWITCH)
   ,.MCAP_EOS_DESIGN_SWITCH(MCAP_EOS_DESIGN_SWITCH)
   ,.MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH(MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH)
   ,.MCAP_GATE_IO_ENABLE_DESIGN_SWITCH(MCAP_GATE_IO_ENABLE_DESIGN_SWITCH)
   ,.SIM_JTAG_IDCODE(SIM_JTAG_IDCODE)
   ,.DEBUG_AXIST_DISABLE_FEATURE_BIT(DEBUG_AXIST_DISABLE_FEATURE_BIT)
   ,.DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS(DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS)
   ,.DEBUG_TL_DISABLE_FC_TIMEOUT(DEBUG_TL_DISABLE_FC_TIMEOUT)
   ,.DEBUG_PL_DISABLE_SCRAMBLING(DEBUG_PL_DISABLE_SCRAMBLING)
   ,.DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL (DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL )
   ,.DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW (DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW )
   ,.DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR(DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR)
   ,.DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR(DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR)
   ,.DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR(DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR)
   ,.DEBUG_PL_SIM_RESET_LFSR(DEBUG_PL_SIM_RESET_LFSR)
   ,.DEBUG_PL_SPARE(DEBUG_PL_SPARE)
   ,.DEBUG_LL_SPARE(DEBUG_LL_SPARE)
   ,.DEBUG_TL_SPARE(DEBUG_TL_SPARE)
   ,.DEBUG_AXI4ST_SPARE(DEBUG_AXI4ST_SPARE)
   ,.DEBUG_CFG_SPARE(DEBUG_CFG_SPARE)
   ,.DEBUG_CAR_SPARE(DEBUG_CAR_SPARE)
   ,.TEST_MODE_PIN_CHAR(TEST_MODE_PIN_CHAR)
   ,.SPARE_BIT0(SPARE_BIT0)
   ,.SPARE_BIT1(SPARE_BIT1)
   ,.SPARE_BIT2(SPARE_BIT2)
   ,.SPARE_BIT3(SPARE_BIT3)
   ,.SPARE_BIT4(SPARE_BIT4)
   ,.SPARE_BIT5(SPARE_BIT5)
   ,.SPARE_BIT6(SPARE_BIT6)
   ,.SPARE_BIT7(SPARE_BIT7)
   ,.SPARE_BIT8(SPARE_BIT8)
   ,.SPARE_BYTE0(SPARE_BYTE0)
   ,.SPARE_BYTE1(SPARE_BYTE1)
   ,.SPARE_BYTE2(SPARE_BYTE2)
   ,.SPARE_BYTE3(SPARE_BYTE3)
   ,.SPARE_WORD0(SPARE_WORD0)
   ,.SPARE_WORD1(SPARE_WORD1)
   ,.SPARE_WORD2(SPARE_WORD2)
   ,.SPARE_WORD3(SPARE_WORD3)

  ) pcie_4_0_pipe_smsw_inst ( 

////////   PIPE Controls ////////////
   .pipe_tx_rcvr_det                   ( pipe_tx0_rcvr_det     ),//(pipe_tx_rcvr_det)
   .pipe_tx_rate                       ( common_commands_out[2:1]   ),//(pipe_tx_rate[1:0])
   .pipe_tx_deemph                     ( common_commands_out[9]     ),//(pipe_tx_deemph)
   .pipe_tx_margin                     ( common_commands_out[6:4]   ),//(pipe_tx_margin[2:0])
   .pipe_tx_swing                      ( common_commands_out[7]     ),//(pipe_tx_swing)
   .pipe_tx_reset                      ( common_commands_out[8]     ),//(pipe_tx_reset)
   .pipe_eq_fs                         ( 6'd40 ),//(pipe_eq_fs[5:0])
   .pipe_eq_lf                         ( 6'd12 ),//(pipe_eq_lf[5:0])

   .pipe_rx_eq_lp_tx_preset (pipe_rx_eq_lp_tx_preset[3:0]),
   .pipe_rx_eq_lp_lf_fs     (pipe_rx_eq_lp_lf_fs[5:0]),
  //-----------------------------
  // PIPE TX BUS Signals[69:0]
  //-----------------------------
  // pipe_tx_0_sigs[69:0]
   .pipe_tx00_data                       ( pipe_tx_0_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx00_char_is_k                  ( pipe_tx_0_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx00_elec_idle                  ( pipe_tx_0_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx00_data_valid                 ( pipe_tx_0_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx00_start_block                ( pipe_tx_0_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx00_sync_header                ( pipe_tx_0_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx00_polarity                   ( pipe_tx_0_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx00_powerdown                  ( pipe_tx_0_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx00_eq_control                 ( pipe_tx00_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_0_sigs[47:44] ),//
   .pipe_tx00_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx00_eq_control                 ( pipe_rx00_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_0_sigs[58:56] ),//
                                       //( pipe_tx_0_sigs[64:59] ),//
                                       //( pipe_tx_0_sigs[68:65] ),//
   .pipe_tx00_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_1_sigs[69:0]
   .pipe_tx01_data                       ( pipe_tx_1_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx01_char_is_k                  ( pipe_tx_1_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx01_elec_idle                  ( pipe_tx_1_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx01_data_valid                 ( pipe_tx_1_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx01_start_block                ( pipe_tx_1_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx01_sync_header                ( pipe_tx_1_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx01_polarity                   ( pipe_tx_1_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx01_powerdown                  ( pipe_tx_1_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx01_eq_control                 ( pipe_tx01_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_1_sigs[47:44] ),//
   .pipe_tx01_eq_deemph                  (  ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx01_eq_control                 ( pipe_rx01_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_1_sigs[58:56] ),//
                                       //( pipe_tx_1_sigs[64:59] ),//
                                       //( pipe_tx_1_sigs[68:65] ),//
   .pipe_tx01_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_2_sigs[69:0]
   .pipe_tx02_data                       ( pipe_tx_2_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx02_char_is_k                  ( pipe_tx_2_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx02_elec_idle                  ( pipe_tx_2_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx02_data_valid                 ( pipe_tx_2_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx02_start_block                ( pipe_tx_2_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx02_sync_header                ( pipe_tx_2_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx02_polarity                   ( pipe_tx_2_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx02_powerdown                  ( pipe_tx_2_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx02_eq_control                 ( pipe_tx02_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_2_sigs[47:44] ),//
   .pipe_tx02_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx02_eq_control                 ( pipe_rx02_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_2_sigs[58:56] ),//
                                       //( pipe_tx_2_sigs[64:59] ),//
                                       //( pipe_tx_2_sigs[68:65] ),//
   .pipe_tx02_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_3_sigs[69:0]
   .pipe_tx03_data                       ( pipe_tx_3_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx03_char_is_k                  ( pipe_tx_3_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx03_elec_idle                  ( pipe_tx_3_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx03_data_valid                 ( pipe_tx_3_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx03_start_block                ( pipe_tx_3_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx03_sync_header                ( pipe_tx_3_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx03_polarity                   ( pipe_tx_3_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx03_powerdown                  ( pipe_tx_3_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx03_eq_control                 ( pipe_tx03_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_3_sigs[47:44] ),//
   .pipe_tx03_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx03_eq_control                 ( pipe_rx03_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_3_sigs[58:56] ),//
                                       //( pipe_tx_3_sigs[64:59] ),//
                                       //( pipe_tx_3_sigs[68:65] ),//
   .pipe_tx03_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_4_sigs[69:0]
   .pipe_tx04_data                       ( pipe_tx_4_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx04_char_is_k                  ( pipe_tx_4_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx04_elec_idle                  ( pipe_tx_4_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx04_data_valid                 ( pipe_tx_4_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx04_start_block                ( pipe_tx_4_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx04_sync_header                ( pipe_tx_4_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx04_polarity                   ( pipe_tx_4_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx04_powerdown                  ( pipe_tx_4_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx04_eq_control                 ( pipe_tx04_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_4_sigs[47:44] ),//
   .pipe_tx04_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx04_eq_control                 ( pipe_rx04_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_4_sigs[58:56] ),//
                                       //( pipe_tx_4_sigs[64:59] ),//
                                       //( pipe_tx_4_sigs[68:65] ),//
   .pipe_tx04_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_5_sigs[69:0]
   .pipe_tx05_data                       ( pipe_tx_5_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx05_char_is_k                  ( pipe_tx_5_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx05_elec_idle                  ( pipe_tx_5_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx05_data_valid                 ( pipe_tx_5_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx05_start_block                ( pipe_tx_5_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx05_sync_header                ( pipe_tx_5_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx05_polarity                   ( pipe_tx_5_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx05_powerdown                  ( pipe_tx_5_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx05_eq_control                 ( pipe_tx05_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_5_sigs[47:44] ),//
   .pipe_tx05_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx05_eq_control                 ( pipe_rx05_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_5_sigs[58:56] ),//
                                       //( pipe_tx_5_sigs[64:59] ),//
                                       //( pipe_tx_5_sigs[68:65] ),//
   .pipe_tx05_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_6_sigs[69:0]
   .pipe_tx06_data                       ( pipe_tx_6_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx06_char_is_k                  ( pipe_tx_6_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx06_elec_idle                  ( pipe_tx_6_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx06_data_valid                 ( pipe_tx_6_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx06_start_block                ( pipe_tx_6_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx06_sync_header                ( pipe_tx_6_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx06_polarity                   ( pipe_tx_6_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx06_powerdown                  ( pipe_tx_6_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx06_eq_control                 ( pipe_tx06_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_6_sigs[47:44] ),//
   .pipe_tx06_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx06_eq_control                 ( pipe_rx06_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_6_sigs[58:56] ),//
                                       //( pipe_tx_6_sigs[64:59] ),//
                                       //( pipe_tx_6_sigs[68:65] ),//
   .pipe_tx06_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_7_sigs[69:0]
   .pipe_tx07_data                       ( pipe_tx_7_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx07_char_is_k                  ( pipe_tx_7_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx07_elec_idle                  ( pipe_tx_7_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx07_data_valid                 ( pipe_tx_7_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx07_start_block                ( pipe_tx_7_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx07_sync_header                ( pipe_tx_7_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx07_polarity                   ( pipe_tx_7_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx07_powerdown                  ( pipe_tx_7_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx07_eq_control                 ( pipe_tx07_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_7_sigs[47:44] ),//
   .pipe_tx07_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx07_eq_control                 ( pipe_rx07_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_7_sigs[58:56] ),//
                                       //( pipe_tx_7_sigs[64:59] ),//
                                       //( pipe_tx_7_sigs[68:65] ),//
   .pipe_tx07_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_8_sigs[69:0]
   .pipe_tx08_data                       ( pipe_tx_8_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx08_char_is_k                  ( pipe_tx_8_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx08_elec_idle                  ( pipe_tx_8_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx08_data_valid                 ( pipe_tx_8_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx08_start_block                ( pipe_tx_8_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx08_sync_header                ( pipe_tx_8_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx08_polarity                   ( pipe_tx_8_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx08_powerdown                  ( pipe_tx_8_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx08_eq_control                 ( pipe_tx08_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_8_sigs[47:44] ),//
   .pipe_tx08_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx08_eq_control                 ( pipe_rx08_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_8_sigs[58:56] ),//
                                       //( pipe_tx_8_sigs[64:59] ),//
                                       //( pipe_tx_8_sigs[68:65] ),//
   .pipe_tx08_compliance                 (  ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_9_sigs[69:0]
   .pipe_tx09_data                       ( pipe_tx_9_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx09_char_is_k                  ( pipe_tx_9_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx09_elec_idle                  ( pipe_tx_9_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx09_data_valid                 ( pipe_tx_9_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx09_start_block                ( pipe_tx_9_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx09_sync_header                ( pipe_tx_9_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx09_polarity                   ( pipe_tx_9_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx09_powerdown                  ( pipe_tx_9_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx09_eq_control                 ( pipe_tx09_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_9_sigs[47:44] ),//
   .pipe_tx09_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx09_eq_control                 ( pipe_rx09_eq_control),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_9_sigs[58:56] ),//
                                       //( pipe_tx_9_sigs[64:59] ),//
                                       //( pipe_tx_9_sigs[68:65] ),//
   .pipe_tx09_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_10_sigs[69:0]
   .pipe_tx10_data                       ( pipe_tx_10_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx10_char_is_k                  ( pipe_tx_10_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx10_elec_idle                  ( pipe_tx_10_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx10_data_valid                 ( pipe_tx_10_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx10_start_block                ( pipe_tx_10_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx10_sync_header                ( pipe_tx_10_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx10_polarity                   ( pipe_tx_10_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx10_powerdown                  ( pipe_tx_10_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx10_eq_control                 ( pipe_tx10_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_10_sigs[47:44] ),//
   .pipe_tx10_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx10_eq_control                 ( pipe_rx10_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_10_sigs[58:56] ),//
                                       //( pipe_tx_10_sigs[64:59] ),//
                                       //( pipe_tx_10_sigs[68:65] ),//
   .pipe_tx10_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_11_sigs[69:0]
   .pipe_tx11_data                       ( pipe_tx_11_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx11_char_is_k                  ( pipe_tx_11_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx11_elec_idle                  ( pipe_tx_11_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx11_data_valid                 ( pipe_tx_11_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx11_start_block                ( pipe_tx_11_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx11_sync_header                ( pipe_tx_11_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx11_polarity                   ( pipe_tx_11_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx11_powerdown                  ( pipe_tx_11_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx11_eq_control                 ( pipe_tx11_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_11_sigs[47:44] ),//
   .pipe_tx11_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx11_eq_control                 ( pipe_rx11_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_11_sigs[58:56] ),//
                                       //( pipe_tx_11_sigs[64:59] ),//
                                       //( pipe_tx_11_sigs[68:65] ),//
   .pipe_tx11_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_12_sigs[69:0]
   .pipe_tx12_data                       ( pipe_tx_12_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx12_char_is_k                  ( pipe_tx_12_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx12_elec_idle                  ( pipe_tx_12_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx12_data_valid                 ( pipe_tx_12_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx12_start_block                ( pipe_tx_12_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx12_sync_header                ( pipe_tx_12_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx12_polarity                   ( pipe_tx_12_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx12_powerdown                  ( pipe_tx_12_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx12_eq_control                 ( pipe_tx12_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_12_sigs[47:44] ),//
   .pipe_tx12_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx12_eq_control                 ( pipe_rx12_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_12_sigs[58:56] ),//
                                       //( pipe_tx_12_sigs[64:59] ),//
                                       //( pipe_tx_12_sigs[68:65] ),//
   .pipe_tx12_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_13_sigs[69:0]
   .pipe_tx13_data                       ( pipe_tx_13_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx13_char_is_k                  ( pipe_tx_13_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx13_elec_idle                  ( pipe_tx_13_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx13_data_valid                 ( pipe_tx_13_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx13_start_block                ( pipe_tx_13_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx13_sync_header                ( pipe_tx_13_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx13_polarity                   ( pipe_tx_13_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx13_powerdown                  ( pipe_tx_13_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx13_eq_control                 ( pipe_tx13_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_13_sigs[47:44] ),//
   .pipe_tx13_eq_deemph                  (  ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx13_eq_control                 ( pipe_rx13_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_13_sigs[58:56] ),//
                                       //( pipe_tx_13_sigs[64:59] ),//
                                       //( pipe_tx_13_sigs[68:65] ),//
   .pipe_tx13_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_14_sigs[69:0]
   .pipe_tx14_data                       ( pipe_tx_14_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx14_char_is_k                  ( pipe_tx_14_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx14_elec_idle                  ( pipe_tx_14_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx14_data_valid                 ( pipe_tx_14_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx14_start_block                ( pipe_tx_14_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx14_sync_header                ( pipe_tx_14_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx14_polarity                   ( pipe_tx_14_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx14_powerdown                  ( pipe_tx_14_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx14_eq_control                 ( pipe_tx14_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_14_sigs[47:44] ),//
   .pipe_tx14_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx14_eq_control                 ( pipe_rx14_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_14_sigs[58:56] ),//
                                       //( pipe_tx_14_sigs[64:59] ),//
                                       //( pipe_tx_14_sigs[68:65] ),//
   .pipe_tx14_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // pipe_tx_15_sigs[69:0]
   .pipe_tx15_data                       ( pipe_tx_15_sigs[31: 0] ),//(pipe_tx00_data[31:0])
   .pipe_tx15_char_is_k                  ( pipe_tx_15_sigs[33:32] ),//(pipe_tx00_char_is_k[1:0])
   .pipe_tx15_elec_idle                  ( pipe_tx_15_sigs[34]    ),//(pipe_tx00_elec_idle)
   .pipe_tx15_data_valid                 ( pipe_tx_15_sigs[35]    ),//(pipe_tx00_data_valid)
   .pipe_tx15_start_block                ( pipe_tx_15_sigs[36]    ),//(pipe_tx00_start_block)
   .pipe_tx15_sync_header                ( pipe_tx_15_sigs[38:37] ),//(pipe_tx00_sync_header[1:0])
   .pipe_rx15_polarity                   ( pipe_tx_15_sigs[39]    ),//(pipe_rx00_polarity)
   .pipe_tx15_powerdown                  ( pipe_tx_15_sigs[41:40] ),//(pipe_tx00_powerdown[1:0])
   .pipe_tx15_eq_control                 ( pipe_tx15_eq_control ),//(pipe_tx00_eq_control[1:0])
                                       //( pipe_tx_15_sigs[47:44] ),//
   .pipe_tx15_eq_deemph                  ( ),//(pipe_tx00_eq_deemph[5:0])
   .pipe_rx15_eq_control                 ( pipe_rx15_eq_control ),//(pipe_rx00_eq_control[1:0])
                                       //( pipe_tx_15_sigs[58:56] ),//
                                       //( pipe_tx_15_sigs[64:59] ),//
                                       //( pipe_tx_15_sigs[68:65] ),//
   .pipe_tx15_compliance                 ( ),//(pipe_tx00_compliance)
  //-----------------------------
  // PIPE RX BUS Signals[83:0]
  //-----------------------------
  // pipe_rx00_sigs[83:0]
   .pipe_rx00_data                         ( pipe_rx_0_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx00_char_is_k                    ( pipe_rx_0_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx00_data_valid                   ( pipe_rx_0_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx00_elec_idle                    ( pipe_rx_0_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx00_start_block                  ( {1'b0, pipe_rx_0_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx00_sync_header                  ( pipe_rx_0_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx00_status                       ( rx_status ),//(pipe_rx00_status[2:0])
   .pipe_rx00_valid                        ( ~pipe_rx_0_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx00_phy_status                   ( phy_status ),//(pipe_rx00_phy_status)
   .pipe_tx00_eq_done                      ( pipe_tx00_eq_done   ),//(pipe_tx00_eq_done)
   .pipe_tx00_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx00_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx00_eq_lp_lf_fs_sel              ( 1'b0    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx00_eq_lp_adapt_done             ( 1'b0   ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx00_eq_done                      ( pipe_rx00_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx01_sigs[83:0]
   .pipe_rx01_data                         ( pipe_rx_1_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx01_char_is_k                    ( pipe_rx_1_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx01_data_valid                   ( pipe_rx_1_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx01_elec_idle                    ( pipe_rx_1_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx01_start_block                  ( {1'b0, pipe_rx_1_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx01_sync_header                  ( pipe_rx_1_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx01_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0  ),//(pipe_rx00_status[2:0])
   .pipe_rx01_valid                        ( ~pipe_rx_1_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx01_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? phy_status : 1'b0  ),//(pipe_rx00_phy_status)
   .pipe_tx01_eq_done                      ( pipe_tx01_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx01_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx01_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx01_eq_lp_lf_fs_sel              ( 1'b0    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx01_eq_lp_adapt_done             ( 1'b0    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx01_eq_done                      ( pipe_rx01_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx02_sigs[83:0]
   .pipe_rx02_data                         ( pipe_rx_2_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx02_char_is_k                    ( pipe_rx_2_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx02_data_valid                   ( pipe_rx_2_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx02_elec_idle                    ( pipe_rx_2_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx02_start_block                  ( {1'b0, pipe_rx_2_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx02_sync_header                  ( pipe_rx_2_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx02_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0  ),//(pipe_rx00_status[2:0])
   .pipe_rx02_valid                        ( ~pipe_rx_2_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx02_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 4 )? phy_status : 1'b0 ),//(pipe_rx00_phy_status)
   .pipe_tx02_eq_done                      ( pipe_tx02_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx02_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx02_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx02_eq_lp_lf_fs_sel              ( 1'b0    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx02_eq_lp_adapt_done             ( 1'b0    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx02_eq_done                      ( pipe_rx02_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx03_sigs[83:0]
   .pipe_rx03_data                         ( pipe_rx_3_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx03_char_is_k                    ( pipe_rx_3_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx03_data_valid                   ( pipe_rx_3_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx03_elec_idle                    ( pipe_rx_3_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx03_start_block                  ( {1'b0, pipe_rx_3_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx03_sync_header                  ( pipe_rx_3_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx03_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0 ),//(pipe_rx00_status[2:0])
   .pipe_rx03_valid                        ( ~pipe_rx_3_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx03_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 4 )? phy_status : 1'b0 ),//(pipe_rx00_phy_status)
   .pipe_tx03_eq_done                      ( pipe_tx03_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx03_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx03_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx03_eq_lp_lf_fs_sel              ( 1'b0    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx03_eq_lp_adapt_done             ( 1'b0    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx03_eq_done                      ( pipe_rx03_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx04_sigs[83:0]
   .pipe_rx04_data                         ( pipe_rx_4_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx04_char_is_k                    ( pipe_rx_4_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx04_data_valid                   ( pipe_rx_4_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx04_elec_idle                    ( pipe_rx_4_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx04_start_block                  ({1'b0,  pipe_rx_4_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx04_sync_header                  ( pipe_rx_4_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx04_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0 ),//(pipe_rx00_status[2:0])
   .pipe_rx04_valid                        ( ~pipe_rx_4_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx04_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 4 )? phy_status : 1'b0    ),//(pipe_rx00_phy_status)
   .pipe_tx04_eq_done                      ( pipe_tx04_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx04_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx04_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx04_eq_lp_lf_fs_sel              ( 1'b0    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx04_eq_lp_adapt_done             ( 1'b0    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx04_eq_done                      ( pipe_rx04_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx05_sigs[83:0]
   .pipe_rx05_data                         ( pipe_rx_5_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx05_char_is_k                    ( pipe_rx_5_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx05_data_valid                   ( pipe_rx_5_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx05_elec_idle                    ( pipe_rx_5_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx05_start_block                  ( {1'b0, pipe_rx_5_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx05_sync_header                  ( pipe_rx_5_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx05_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0 ),//(pipe_rx00_status[2:0])
   .pipe_rx05_valid                        ( ~pipe_rx_5_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx05_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 4 )? phy_status : 1'b0    ),//(pipe_rx00_phy_status)
   .pipe_tx05_eq_done                      ( pipe_tx05_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx05_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx05_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx05_eq_lp_lf_fs_sel              ( 1'b0    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx05_eq_lp_adapt_done             ( 1'b0    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx05_eq_done                      ( pipe_rx05_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx06_sigs[83:0]
   .pipe_rx06_data                         ( pipe_rx_6_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx06_char_is_k                    ( pipe_rx_6_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx06_data_valid                   ( pipe_rx_6_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx06_elec_idle                    ( pipe_rx_6_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx06_start_block                  ( {1'b0, pipe_rx_6_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx06_sync_header                  ( pipe_rx_6_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx06_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0 ),//(pipe_rx00_status[2:0])
   .pipe_rx06_valid                        ( ~pipe_rx_6_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx06_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 4 )? phy_status : 1'b0    ),//(pipe_rx00_phy_status)
   .pipe_tx06_eq_done                      ( pipe_tx06_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx06_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx06_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx06_eq_lp_lf_fs_sel              ( 1'b1    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx06_eq_lp_adapt_done             ( 1'b1    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx06_eq_done                      ( pipe_rx06_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx07_sigs[83:0]
   .pipe_rx07_data                         ( pipe_rx_7_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx07_char_is_k                    ( pipe_rx_7_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx07_data_valid                   ( pipe_rx_7_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx07_elec_idle                    ( pipe_rx_7_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx07_start_block                  ( {1'b0, pipe_rx_7_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx07_sync_header                  ( pipe_rx_7_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx07_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0 ),//(pipe_rx00_status[2:0])
   .pipe_rx07_valid                        ( ~pipe_rx_7_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx07_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 4 )? phy_status : 1'b0     ),//(pipe_rx00_phy_status)
   .pipe_tx07_eq_done                      ( pipe_tx07_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx07_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx07_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx07_eq_lp_lf_fs_sel              ( 1'b1   ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx07_eq_lp_adapt_done             ( 1'b1    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx07_eq_done                      ( pipe_rx07_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx08_sigs[83:0]
   .pipe_rx08_data                         ( pipe_rx_8_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx08_char_is_k                    ( pipe_rx_8_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx08_data_valid                   ( pipe_rx_8_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx08_elec_idle                    ( pipe_rx_8_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx08_start_block                  ( {1'b0, pipe_rx_8_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx08_sync_header                  ( pipe_rx_8_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx08_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0 ),//(pipe_rx00_status[2:0])
   .pipe_rx08_valid                        ( ~pipe_rx_8_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx08_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 8 )? phy_status : 1'b0  ),//(pipe_rx00_phy_status)
   .pipe_tx08_eq_done                      ( pipe_tx08_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx08_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx08_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx08_eq_lp_lf_fs_sel              ( 1'b1    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx08_eq_lp_adapt_done             ( 1'b1    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx08_eq_done                      ( pipe_rx08_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx09_sigs[83:0]
   .pipe_rx09_data                         ( pipe_rx_9_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx09_char_is_k                    ( pipe_rx_9_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx09_data_valid                   ( pipe_rx_9_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx09_elec_idle                    ( pipe_rx_9_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx09_start_block                  ( {1'b0, pipe_rx_9_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx09_sync_header                  ( pipe_rx_9_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx09_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0  ),//(pipe_rx00_status[2:0])
   .pipe_rx09_valid                        ( ~pipe_rx_9_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx09_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 8 )? phy_status : 1'b0    ),//(pipe_rx00_phy_status)
   .pipe_tx09_eq_done                      ( pipe_tx09_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx09_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx09_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx09_eq_lp_lf_fs_sel              ( 1'b1    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx09_eq_lp_adapt_done             ( 1'b1    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx09_eq_done                      ( pipe_rx09_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx10_sigs[83:0]
   .pipe_rx10_data                         ( pipe_rx_10_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx10_char_is_k                    ( pipe_rx_10_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx10_data_valid                   ( pipe_rx_10_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx10_elec_idle                    ( pipe_rx_10_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx10_start_block                  ( {1'b0, pipe_rx_10_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx10_sync_header                  ( pipe_rx_10_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx10_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0 ),//(pipe_rx00_status[2:0])
   .pipe_rx10_valid                        ( ~pipe_rx_10_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx10_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 8 )? phy_status : 1'b0   ),//(pipe_rx00_phy_status)
   .pipe_tx10_eq_done                      ( pipe_tx10_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx10_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx10_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx10_eq_lp_lf_fs_sel              ( 1'b1    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx10_eq_lp_adapt_done             ( 1'b1    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx10_eq_done                      ( pipe_rx10_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx11_sigs[83:0]
   .pipe_rx11_data                         ( pipe_rx_11_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx11_char_is_k                    ( pipe_rx_11_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx11_data_valid                   ( pipe_rx_11_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx11_elec_idle                    ( pipe_rx_11_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx11_start_block                  ( {1'b0, pipe_rx_11_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx11_sync_header                  ( pipe_rx_11_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx11_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0 ),//(pipe_rx00_status[2:0])
   .pipe_rx11_valid                        ( ~pipe_rx_11_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx11_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 8 )? phy_status : 1'b0    ),//(pipe_rx00_phy_status)
   .pipe_tx11_eq_done                      ( pipe_tx11_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx11_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx11_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx11_eq_lp_lf_fs_sel              ( 1'b1    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx11_eq_lp_adapt_done             ( 1'b1    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx11_eq_done                      ( pipe_rx11_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx12_sigs[83:0]
   .pipe_rx12_data                         ( pipe_rx_12_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx12_char_is_k                    ( pipe_rx_12_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx12_data_valid                   ( pipe_rx_12_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx12_elec_idle                    ( pipe_rx_12_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx12_start_block                  ( {1'b0, pipe_rx_12_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx12_sync_header                  ( pipe_rx_12_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx12_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0 ),//(pipe_rx00_status[2:0])
   .pipe_rx12_valid                        ( ~pipe_rx_12_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx12_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 8 )? phy_status : 1'b0    ),//(pipe_rx00_phy_status)
   .pipe_tx12_eq_done                      ( pipe_tx12_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx12_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx12_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx12_eq_lp_lf_fs_sel              ( 1'b1    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx12_eq_lp_adapt_done             ( 1'b1    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx12_eq_done                      ( pipe_rx12_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx13_sigs[83:0]
   .pipe_rx13_data                         ( pipe_rx_13_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx13_char_is_k                    ( pipe_rx_13_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx13_data_valid                   ( pipe_rx_13_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx13_elec_idle                    ( pipe_rx_13_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx13_start_block                  ( {1'b0, pipe_rx_13_sigs[36]}    ),//(pipe_rx00_start_block[1:0])
   .pipe_rx13_sync_header                  ( pipe_rx_13_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx13_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0 ),//(pipe_rx00_status[2:0])
   .pipe_rx13_valid                        ( ~pipe_rx_13_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx13_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 8 )? phy_status : 1'b0    ),//(pipe_rx00_phy_status)
   .pipe_tx13_eq_done                      ( pipe_tx13_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx13_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx13_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx13_eq_lp_lf_fs_sel              ( 1'b1    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx13_eq_lp_adapt_done             ( 1'b1    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx13_eq_done                      ( pipe_rx13_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx14_sigs[83:0]
   .pipe_rx14_data                         ( pipe_rx_14_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx14_char_is_k                    ( pipe_rx_14_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx14_data_valid                   ( pipe_rx_14_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx14_elec_idle                    ( pipe_rx_14_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx14_start_block                  ( {1'b0, pipe_rx_14_sigs[36] }   ),//(pipe_rx00_start_block[1:0])
   .pipe_rx14_sync_header                  ( pipe_rx_14_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx14_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0 ),//(pipe_rx00_status[2:0])
   .pipe_rx14_valid                        ( ~pipe_rx_14_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx14_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 8 )? phy_status : 1'b0     ),//(pipe_rx00_phy_status)
   .pipe_tx14_eq_done                      ( pipe_tx14_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx14_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx14_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx14_eq_lp_lf_fs_sel              ( 1'b1    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx14_eq_lp_adapt_done             ( 1'b1    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx14_eq_done                      ( pipe_rx14_eq_done    ),//(pipe_rx00_eq_done)
  //-----------------------------
  // pipe_rx15_sigs[83:0]
   .pipe_rx15_data                         ( pipe_rx_15_sigs[31: 0] ),//(pipe_rx00_data[31:0])
   .pipe_rx15_char_is_k                    ( pipe_rx_15_sigs[33:32] ),//(pipe_rx00_char_is_k[1:0])
   .pipe_rx15_data_valid                   ( pipe_rx_15_sigs[35]    ),//(pipe_rx00_data_valid)
   .pipe_rx15_elec_idle                    ( pipe_rx_15_sigs[34]    ),//(pipe_rx00_elec_idle)
   .pipe_rx15_start_block                  ( {1'b0, pipe_rx_15_sigs[36] }   ),//(pipe_rx00_start_block[1:0])
   .pipe_rx15_sync_header                  ( pipe_rx_15_sigs[38:37] ),//(pipe_rx00_sync_header[1:0])
   .pipe_rx15_status                       ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 2 )? rx_status : 3'b0 ),//(pipe_rx00_status[2:0])
   .pipe_rx15_valid                        ( ~pipe_rx_15_sigs[34]    ),//(pipe_rx00_valid)
   .pipe_rx15_phy_status                   ( (PL_LINK_CAP_MAX_LINK_WIDTH >= 8 )? phy_status : 1'b0    ),//(pipe_rx00_phy_status)
   .pipe_tx15_eq_done                      ( pipe_tx15_eq_done    ),//(pipe_tx00_eq_done)
   .pipe_tx15_eq_coeff                     ( 18'h00904 ),//(pipe_tx00_eq_coeff[17:0])
   .pipe_rx15_eq_lp_new_tx_coeff_or_preset ( 18'h05 ),//(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   .pipe_rx15_eq_lp_lf_fs_sel              ( 1'b1    ),//(pipe_rx00_eq_lp_lf_fs_sel)
   .pipe_rx15_eq_lp_adapt_done             ( 1'b1    ),//(pipe_rx00_eq_lp_adapt_done)
   .pipe_rx15_eq_done                      ( pipe_rx15_eq_done    )//(pipe_rx00_eq_done)

   //,.pipe_rx08_data( pipe_tx_rate==2'b11 ? pipe_rx00_data[63:32] : pipe_rx08_data[31:0] )
   //,.pipe_rx09_data( pipe_tx_rate==2'b11 ? pipe_rx01_data[63:32] : pipe_rx09_data[31:0] )
   //,.pipe_rx10_data( pipe_tx_rate==2'b11 ? pipe_rx02_data[63:32] : pipe_rx10_data[31:0] )
   //,.pipe_rx11_data( pipe_tx_rate==2'b11 ? pipe_rx03_data[63:32] : pipe_rx11_data[31:0] )
   //,.pipe_rx12_data( pipe_tx_rate==2'b11 ? pipe_rx04_data[63:32] : pipe_rx12_data[31:0] )
   //,.pipe_rx13_data( pipe_tx_rate==2'b11 ? pipe_rx05_data[63:32] : pipe_rx13_data[31:0] )
   //,.pipe_rx14_data( pipe_tx_rate==2'b11 ? pipe_rx06_data[63:32] : pipe_rx14_data[31:0] )
   //,.pipe_rx15_data( pipe_tx_rate==2'b11 ? pipe_rx07_data[63:32] : pipe_rx15_data[31:0] )
   // -------------------------------------------------------------------------------------
   ,.pl_gen2_upstream_prefer_deemph(pl_gen2_upstream_prefer_deemph)
   ,.pl_eq_in_progress(pl_eq_in_progress)
   ,.pl_eq_phase(pl_eq_phase[1:0])
   ,.pl_eq_reset_eieos_count(1'b0)
   ,.pl_redo_eq(pl_redo_eq)
   ,.pl_redo_eq_speed(pl_redo_eq_speed)
   ,.pl_eq_mismatch(pl_eq_mismatch)
   ,.pl_redo_eq_pending(pl_redo_eq_pending)
   ,.m_axis_cq_tdata(m_axis_cq_tdata[AXI4_DATA_WIDTH-1:0])
   ,.s_axis_cc_tdata(s_axis_cc_tdata[AXI4_DATA_WIDTH-1:0])
   ,.s_axis_rq_tdata(s_axis_rq_tdata[AXI4_DATA_WIDTH-1:0])
   ,.m_axis_rc_tdata(m_axis_rc_tdata[AXI4_DATA_WIDTH-1:0])
   ,.m_axis_cq_tuser(m_axis_cq_tuser[AXI4_CQ_TUSER_WIDTH-1:0])
   ,.s_axis_cc_tuser(s_axis_cc_tuser[AXI4_CC_TUSER_WIDTH-1:0])
   ,.m_axis_cq_tlast(m_axis_cq_tlast)
   ,.s_axis_rq_tlast(s_axis_rq_tlast)
   ,.m_axis_rc_tlast(m_axis_rc_tlast)
   ,.s_axis_cc_tlast(s_axis_cc_tlast)
   ,.pcie_cq_np_req(pcie_cq_np_req[1:0])
   ,.pcie_cq_np_req_count(pcie_cq_np_req_count[5:0])
   ,.s_axis_rq_tuser(s_axis_rq_tuser[AXI4_RQ_TUSER_WIDTH-1:0])
   ,.m_axis_rc_tuser(m_axis_rc_tuser[AXI4_RC_TUSER_WIDTH-1:0])
   ,.m_axis_cq_tkeep(m_axis_cq_tkeep[AXI4_TKEEP_WIDTH-1:0])
   ,.s_axis_cc_tkeep(s_axis_cc_tkeep[AXI4_TKEEP_WIDTH-1:0])
   ,.s_axis_rq_tkeep(s_axis_rq_tkeep[AXI4_TKEEP_WIDTH-1:0])
   ,.m_axis_rc_tkeep(m_axis_rc_tkeep[AXI4_TKEEP_WIDTH-1:0])
   ,.m_axis_cq_tvalid(m_axis_cq_tvalid)
   ,.s_axis_cc_tvalid(s_axis_cc_tvalid)
   ,.s_axis_rq_tvalid(s_axis_rq_tvalid)
   ,.m_axis_rc_tvalid(m_axis_rc_tvalid)
   ,.m_axis_cq_tready({AXI4_CQ_TREADY_WIDTH{m_axis_cq_tready}})
   ,.s_axis_cc_tready(s_axis_cc_tready)
   ,.s_axis_rq_tready(s_axis_rq_tready)
   ,.m_axis_rc_tready({AXI4_RC_TREADY_WIDTH{m_axis_rc_tready}})
   ,.pcie_rq_seq_num0(pcie_rq_seq_num0[5:0])
   ,.pcie_rq_seq_num_vld0(pcie_rq_seq_num_vld0)
   ,.pcie_rq_seq_num1(pcie_rq_seq_num1[5:0])
   ,.pcie_rq_seq_num_vld1(pcie_rq_seq_num_vld1)
   ,.pcie_rq_tag0(pcie_rq_tag0[7:0])
   ,.pcie_rq_tag_vld0(pcie_rq_tag_vld0)
   ,.pcie_rq_tag1(pcie_rq_tag1[7:0])
   ,.pcie_rq_tag_vld1(pcie_rq_tag_vld1)
   ,.pcie_tfc_nph_av(pcie_tfc_nph_av[3:0])
   ,.pcie_tfc_npd_av(pcie_tfc_npd_av[3:0])
   ,.pcie_rq_tag_av(pcie_rq_tag_av[3:0])
   ,.axi_user_out( )
   ,.axi_user_in(8'h00)
   ,.cfg_mgmt_addr(cfg_mgmt_addr[9:0])
   ,.cfg_mgmt_function_number(cfg_mgmt_function_number[7:0])
   ,.cfg_mgmt_write(cfg_mgmt_write)
   ,.cfg_mgmt_write_data(cfg_mgmt_write_data[31:0])
   ,.cfg_mgmt_byte_enable(cfg_mgmt_byte_enable[3:0])
   ,.cfg_mgmt_read(cfg_mgmt_read)
   ,.cfg_mgmt_read_data(cfg_mgmt_read_data[31:0])
   ,.cfg_mgmt_read_write_done(cfg_mgmt_read_write_done)
   ,.cfg_mgmt_debug_access(cfg_mgmt_debug_access)
   ,.cfg_phy_link_down(cfg_phy_link_down)
   ,.cfg_phy_link_status(cfg_phy_link_status[1:0])
   ,.cfg_negotiated_width(cfg_negotiated_width[2:0])
   ,.cfg_current_speed(cfg_current_speed[1:0])
   ,.cfg_max_payload(cfg_max_payload[1:0])
   ,.cfg_max_read_req(cfg_max_read_req[2:0])
   ,.cfg_function_status(cfg_function_status[15:0])
   ,.cfg_function_power_state(cfg_function_power_state[11:0])
   ,.cfg_link_power_state(cfg_link_power_state[1:0])
   ,.cfg_err_cor_out(cfg_err_cor_out)
   ,.cfg_err_nonfatal_out(cfg_err_nonfatal_out)
   ,.cfg_err_fatal_out(cfg_err_fatal_out)
   ,.cfg_local_error_valid(cfg_local_error_valid)
   ,.cfg_local_error_out(cfg_local_error_out[4:0])
   ,.cfg_ltr_enable()
   ,.cfg_ltssm_state(cfg_ltssm_state[5:0])
   ,.cfg_rx_pm_state(cfg_rx_pm_state[1:0])
   ,.cfg_tx_pm_state(cfg_tx_pm_state[1:0])
   ,.cfg_rcb_status(cfg_rcb_status[3:0])
   ,.cfg_obff_enable(cfg_obff_enable[1:0])
   ,.cfg_pl_status_change(cfg_pl_status_change)
   ,.cfg_tph_requester_enable(cfg_tph_requester_enable[3:0])
   ,.cfg_tph_st_mode(cfg_tph_st_mode[11:0])
   ,.cfg_msg_received(cfg_msg_received)
   ,.cfg_msg_received_data(cfg_msg_received_data[7:0])
   ,.cfg_msg_received_type(cfg_msg_received_type[4:0])
   ,.cfg_msg_transmit(cfg_msg_transmit_int)
   ,.cfg_msg_transmit_type(cfg_msg_transmit_type[2:0])
   ,.cfg_msg_transmit_data(cfg_msg_transmit_data[31:0])
   ,.cfg_msg_transmit_done(cfg_msg_transmit_done)
   ,.cfg_fc_ph(cfg_fc_ph[7:0])
   ,.cfg_fc_pd(cfg_fc_pd[11:0])
   ,.cfg_fc_nph(cfg_fc_nph[7:0])
   ,.cfg_fc_npd(cfg_fc_npd[11:0])
   ,.cfg_fc_cplh(cfg_fc_cplh[7:0])
   ,.cfg_fc_cpld(cfg_fc_cpld[11:0])
   ,.cfg_fc_sel(cfg_fc_sel[2:0])
   ,.cfg_hot_reset_in(cfg_hot_reset_in)
   ,.cfg_hot_reset_out(cfg_hot_reset_out)
   ,.cfg_config_space_enable(cfg_config_space_enable)
   ,.cfg_dsn(cfg_dsn[63:0])
   ,.cfg_dev_id_pf0(cfg_dev_id_pf0[15:0])
   ,.cfg_dev_id_pf1(cfg_dev_id_pf1[15:0])
   ,.cfg_dev_id_pf2(cfg_dev_id_pf2[15:0])
   ,.cfg_dev_id_pf3(cfg_dev_id_pf3[15:0])
   ,.cfg_vend_id(cfg_vend_id[15:0])
   ,.cfg_rev_id_pf0(cfg_rev_id_pf0[7:0])
   ,.cfg_rev_id_pf1(cfg_rev_id_pf1[7:0])
   ,.cfg_rev_id_pf2(cfg_rev_id_pf2[7:0])
   ,.cfg_rev_id_pf3(cfg_rev_id_pf3[7:0])
   ,.cfg_subsys_id_pf0(cfg_subsys_id_pf0[15:0])
   ,.cfg_subsys_id_pf1(cfg_subsys_id_pf1[15:0])
   ,.cfg_subsys_id_pf2(cfg_subsys_id_pf2[15:0])
   ,.cfg_subsys_id_pf3(cfg_subsys_id_pf3[15:0])
   ,.cfg_subsys_vend_id(cfg_subsys_vend_id[15:0])
   ,.cfg_ds_port_number(cfg_ds_port_number[7:0])
   ,.cfg_ds_bus_number(cfg_ds_bus_number[7:0])
   ,.cfg_ds_device_number(cfg_ds_device_number[4:0])
   ,.cfg_ds_function_number(3'b0)
   ,.cfg_bus_number(cfg_bus_number[7:0])
   ,.cfg_power_state_change_ack(cfg_power_state_change_ack)
   ,.cfg_power_state_change_interrupt(cfg_power_state_change_interrupt)
   ,.cfg_err_cor_in(cfg_err_cor_in)
   ,.cfg_err_uncor_in(cfg_err_uncor_in)
   ,.cfg_flr_done(cfg_flr_done[3:0])
   ,.cfg_vf_flr_in_process(cfg_vf_flr_in_process[251:0])   
   ,.cfg_vf_flr_done(cfg_vf_flr_done)                      
   ,.cfg_vf_flr_func_num(cfg_vf_flr_func_num[7:0])
   ,.cfg_vf_status(cfg_vf_status[503:0])                   
   ,.cfg_vf_power_state(cfg_vf_power_state[755:0])         
   ,.cfg_vf_tph_requester_enable( cfg_vf_tph_requester_enable[251:0])
   ,.cfg_vf_tph_st_mode(cfg_vf_tph_st_mode[755:0])         
   ,.cfg_interrupt_msix_vf_enable(cfg_interrupt_msix_vf_enable[251:0])
   ,.cfg_interrupt_msix_vf_mask(cfg_interrupt_msix_vf_mask[251:0])
   ,.cfg_flr_in_process(cfg_flr_in_process[3:0])
   ,.cfg_req_pm_transition_l23_ready(cfg_req_pm_transition_l23_ready)
   ,.cfg_link_training_enable(cfg_link_training_enable)
   ,.cfg_interrupt_int(cfg_interrupt_int[3:0])
   ,.cfg_interrupt_sent(cfg_interrupt_sent)
   ,.cfg_interrupt_pending(cfg_interrupt_pending[3:0])
   ,.cfg_interrupt_msi_enable(cfg_interrupt_msi_enable[3:0])
   ,.cfg_interrupt_msi_int(cfg_interrupt_msi_int[31:0])
   ,.cfg_interrupt_msi_sent(cfg_interrupt_msi_sent)
   ,.cfg_interrupt_msi_fail(cfg_interrupt_msi_fail)
   ,.cfg_interrupt_msi_mmenable(cfg_interrupt_msi_mmenable[11:0])
   ,.cfg_interrupt_msi_pending_status(cfg_interrupt_msi_pending_status[31:0])
   ,.cfg_interrupt_msi_pending_status_function_num(cfg_interrupt_msi_pending_status_function_num[1:0])
   ,.cfg_interrupt_msi_pending_status_data_enable(cfg_interrupt_msi_pending_status_data_enable)
   ,.cfg_interrupt_msi_mask_update(cfg_interrupt_msi_mask_update)
   ,.cfg_interrupt_msi_select(cfg_interrupt_msi_select[1:0])
   ,.cfg_interrupt_msi_data(cfg_interrupt_msi_data[31:0])
   ,.cfg_interrupt_msix_enable(cfg_interrupt_msix_enable[3:0])
   ,.cfg_interrupt_msix_mask(cfg_interrupt_msix_mask[3:0])
   ,.cfg_interrupt_msix_address(cfg_interrupt_msix_address[63:0])
   ,.cfg_interrupt_msix_data(cfg_interrupt_msix_data[31:0])
   ,.cfg_interrupt_msix_int(cfg_interrupt_msix_int)
   ,.cfg_interrupt_msix_vec_pending(cfg_interrupt_msix_vec_pending[1:0])
   ,.cfg_interrupt_msix_vec_pending_status(cfg_interrupt_msix_vec_pending_status)
   ,.cfg_interrupt_msi_attr(cfg_interrupt_msi_attr[2:0])
   ,.cfg_interrupt_msi_tph_present(cfg_interrupt_msi_tph_present)
   ,.cfg_interrupt_msi_tph_type(cfg_interrupt_msi_tph_type[1:0])
   ,.cfg_interrupt_msi_tph_st_tag(cfg_interrupt_msi_tph_st_tag[7:0])
   ,.cfg_interrupt_msi_function_number(cfg_interrupt_msi_function_number[7:0])
   ,.cfg_ext_read_received(cfg_ext_read_received)
   ,.cfg_ext_write_received(cfg_ext_write_received)
   ,.cfg_ext_register_number(cfg_ext_register_number[9:0])
   ,.cfg_ext_function_number(cfg_ext_function_number[7:0])
   ,.cfg_ext_write_data(cfg_ext_write_data[31:0])
   ,.cfg_ext_write_byte_enable(cfg_ext_write_byte_enable[3:0])
   ,.cfg_ext_read_data(cfg_ext_read_data[31:0])
   ,.cfg_ext_read_data_valid(cfg_ext_read_data_valid)
   ,.cfg_pm_aspm_l1_entry_reject(cfg_pm_aspm_l1_entry_reject)
   ,.cfg_pm_aspm_tx_l0s_entry_disable(cfg_pm_aspm_tx_l0s_entry_disable)
   ,.user_tph_stt_func_num(8'h00)
   ,.user_tph_stt_index(6'b0)
   ,.user_tph_stt_rd_en(1'b0)
   ,.user_tph_stt_rd_data()
   ,.conf_req_type(conf_req_type[1:0])
   ,.conf_req_reg_num(conf_req_reg_num[3:0])
   ,.conf_req_data(conf_req_data[31:0])
   ,.conf_req_valid(conf_req_valid)
   ,.conf_req_ready(conf_req_ready)
   ,.conf_resp_rdata(conf_resp_rdata[31:0])
   ,.conf_resp_valid(conf_resp_valid)
   ,.conf_mcap_design_switch(conf_mcap_design_switch)
   ,.conf_mcap_eos(conf_mcap_eos)
   ,.conf_mcap_in_use_by_pcie(conf_mcap_in_use_by_pcie)
   ,.conf_mcap_request_by_conf(conf_mcap_request_by_conf)

   ,.drp_clk('h0)
   ,.drp_en('h0)
   ,.drp_we('h0)
   ,.drp_addr('h0)
   ,.drp_di('h0)
   ,.drp_rdy()
   ,.drp_do()

   ,.pipe_clk(pipe_clk)
   ,.core_clk(core_clk)
   ,.user_clk(user_clk)
   ,.user_clk2(user_clk2)
   ,.user_clk_en(user_clk_en)
   ,.mcap_clk(mcap_clk)
   ,.mcap_rst_b(mcap_rst_b)
   ,.pcie_perst0_b(pcie_perst0_b)
   ,.pcie_perst1_b(pcie_perst1_b)
   ,.phy_rdy(phy_rdy)

  );
  
  reg [3:0] pipe_rx00_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx01_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx02_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx03_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx04_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx05_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx06_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx07_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx08_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx09_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx10_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx11_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx12_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx13_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx14_eq_control_reg = 4'b0;
  reg [3:0] pipe_rx15_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx00_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx01_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx02_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx03_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx04_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx05_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx06_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx07_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx08_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx09_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx10_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx11_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx12_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx13_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx14_eq_control_reg = 4'b0;
  reg [3:0] pipe_tx15_eq_control_reg = 4'b0;

  always @ (posedge pipe_clk)
  begin
   pipe_rx00_eq_control_reg     <= {pipe_rx00_eq_control_reg[1:0], pipe_rx00_eq_control};
   pipe_rx01_eq_control_reg     <= {pipe_rx01_eq_control_reg[1:0], pipe_rx01_eq_control};
   pipe_rx02_eq_control_reg     <= {pipe_rx02_eq_control_reg[1:0], pipe_rx02_eq_control};
   pipe_rx03_eq_control_reg     <= {pipe_rx03_eq_control_reg[1:0], pipe_rx03_eq_control};
   pipe_rx04_eq_control_reg     <= {pipe_rx04_eq_control_reg[1:0], pipe_rx04_eq_control};
   pipe_rx05_eq_control_reg     <= {pipe_rx05_eq_control_reg[1:0], pipe_rx05_eq_control};
   pipe_rx06_eq_control_reg     <= {pipe_rx06_eq_control_reg[1:0], pipe_rx06_eq_control};
   pipe_rx07_eq_control_reg     <= {pipe_rx07_eq_control_reg[1:0], pipe_rx07_eq_control};
   pipe_rx08_eq_control_reg     <= {pipe_rx08_eq_control_reg[1:0], pipe_rx08_eq_control};
   pipe_rx09_eq_control_reg     <= {pipe_rx09_eq_control_reg[1:0], pipe_rx09_eq_control};
   pipe_rx10_eq_control_reg     <= {pipe_rx10_eq_control_reg[1:0], pipe_rx10_eq_control};
   pipe_rx11_eq_control_reg     <= {pipe_rx11_eq_control_reg[1:0], pipe_rx11_eq_control};
   pipe_rx12_eq_control_reg     <= {pipe_rx12_eq_control_reg[1:0], pipe_rx12_eq_control};
   pipe_rx13_eq_control_reg     <= {pipe_rx13_eq_control_reg[1:0], pipe_rx13_eq_control};
   pipe_rx14_eq_control_reg     <= {pipe_rx14_eq_control_reg[1:0], pipe_rx14_eq_control};
   pipe_rx15_eq_control_reg     <= {pipe_rx15_eq_control_reg[1:0], pipe_rx15_eq_control};

   pipe_tx00_eq_control_reg     <= {pipe_tx00_eq_control_reg[1:0], pipe_tx00_eq_control};
   pipe_tx01_eq_control_reg     <= {pipe_tx01_eq_control_reg[1:0], pipe_tx01_eq_control};
   pipe_tx02_eq_control_reg     <= {pipe_tx02_eq_control_reg[1:0], pipe_tx02_eq_control};
   pipe_tx03_eq_control_reg     <= {pipe_tx03_eq_control_reg[1:0], pipe_tx03_eq_control};
   pipe_tx04_eq_control_reg     <= {pipe_tx04_eq_control_reg[1:0], pipe_tx04_eq_control};
   pipe_tx05_eq_control_reg     <= {pipe_tx05_eq_control_reg[1:0], pipe_tx05_eq_control};
   pipe_tx06_eq_control_reg     <= {pipe_tx06_eq_control_reg[1:0], pipe_tx06_eq_control};
   pipe_tx07_eq_control_reg     <= {pipe_tx07_eq_control_reg[1:0], pipe_tx07_eq_control};
   pipe_tx08_eq_control_reg     <= {pipe_tx08_eq_control_reg[1:0], pipe_tx08_eq_control};
   pipe_tx09_eq_control_reg     <= {pipe_tx09_eq_control_reg[1:0], pipe_tx09_eq_control};
   pipe_tx10_eq_control_reg     <= {pipe_tx10_eq_control_reg[1:0], pipe_tx10_eq_control};
   pipe_tx11_eq_control_reg     <= {pipe_tx11_eq_control_reg[1:0], pipe_tx11_eq_control};
   pipe_tx12_eq_control_reg     <= {pipe_tx12_eq_control_reg[1:0], pipe_tx12_eq_control};
   pipe_tx13_eq_control_reg     <= {pipe_tx13_eq_control_reg[1:0], pipe_tx13_eq_control};
   pipe_tx14_eq_control_reg     <= {pipe_tx14_eq_control_reg[1:0], pipe_tx14_eq_control};
   pipe_tx15_eq_control_reg     <= {pipe_tx15_eq_control_reg[1:0], pipe_tx15_eq_control};

  end
  
  
  // generate rx*_eq_done
  assign pipe_rx00_eq_done = (pipe_rx00_eq_control_reg[3:2] != pipe_rx00_eq_control)? 1'b1 : 1'b0;
  assign pipe_rx01_eq_done = (pipe_rx01_eq_control_reg[3:2] != pipe_rx01_eq_control)? 1'b1 : 1'b0;
  assign pipe_rx02_eq_done = (pipe_rx02_eq_control_reg[3:2] != pipe_rx02_eq_control)? 1'b1 : 1'b0;
  assign pipe_rx03_eq_done = (pipe_rx03_eq_control_reg[3:2] != pipe_rx03_eq_control)? 1'b1 : 1'b0;
  assign pipe_rx04_eq_done = (pipe_rx04_eq_control_reg[3:2] != pipe_rx04_eq_control)? 1'b1 : 1'b0;
  assign pipe_rx05_eq_done = (pipe_rx05_eq_control_reg[3:2] != pipe_rx05_eq_control)? 1'b1 : 1'b0;
  assign pipe_rx06_eq_done = (pipe_rx06_eq_control_reg[3:2] != pipe_rx06_eq_control)? 1'b1 : 1'b0;
  assign pipe_rx07_eq_done = (pipe_rx07_eq_control_reg[3:2] != pipe_rx07_eq_control)? 1'b1 : 1'b0; 
  assign pipe_rx08_eq_done = (pipe_rx08_eq_control_reg[3:2] != pipe_rx08_eq_control)? 1'b1 : 1'b0; 
  assign pipe_rx09_eq_done = (pipe_rx09_eq_control_reg[3:2] != pipe_rx09_eq_control)? 1'b1 : 1'b0; 
  assign pipe_rx10_eq_done = (pipe_rx10_eq_control_reg[3:2] != pipe_rx10_eq_control)? 1'b1 : 1'b0; 
  assign pipe_rx11_eq_done = (pipe_rx11_eq_control_reg[3:2] != pipe_rx11_eq_control)? 1'b1 : 1'b0; 
  assign pipe_rx12_eq_done = (pipe_rx12_eq_control_reg[3:2] != pipe_rx12_eq_control)? 1'b1 : 1'b0; 
  assign pipe_rx13_eq_done = (pipe_rx13_eq_control_reg[3:2] != pipe_rx13_eq_control)? 1'b1 : 1'b0; 
  assign pipe_rx14_eq_done = (pipe_rx14_eq_control_reg[3:2] != pipe_rx14_eq_control)? 1'b1 : 1'b0; 
  assign pipe_rx15_eq_done = (pipe_rx15_eq_control_reg[3:2] != pipe_rx15_eq_control)? 1'b1 : 1'b0; 
  // generate tx*_eq_done
  assign pipe_tx00_eq_done = (pipe_tx00_eq_control_reg[3:2] != pipe_tx00_eq_control)? 1'b1 : 1'b0;
  assign pipe_tx01_eq_done = (pipe_tx01_eq_control_reg[3:2] != pipe_tx01_eq_control)? 1'b1 : 1'b0;
  assign pipe_tx02_eq_done = (pipe_tx02_eq_control_reg[3:2] != pipe_tx02_eq_control)? 1'b1 : 1'b0;
  assign pipe_tx03_eq_done = (pipe_tx03_eq_control_reg[3:2] != pipe_tx03_eq_control)? 1'b1 : 1'b0;
  assign pipe_tx04_eq_done = (pipe_tx04_eq_control_reg[3:2] != pipe_tx04_eq_control)? 1'b1 : 1'b0;
  assign pipe_tx05_eq_done = (pipe_tx05_eq_control_reg[3:2] != pipe_tx05_eq_control)? 1'b1 : 1'b0;
  assign pipe_tx06_eq_done = (pipe_tx06_eq_control_reg[3:2] != pipe_tx06_eq_control)? 1'b1 : 1'b0;
  assign pipe_tx07_eq_done = (pipe_tx07_eq_control_reg[3:2] != pipe_tx07_eq_control)? 1'b1 : 1'b0; 
  assign pipe_tx08_eq_done = (pipe_tx08_eq_control_reg[3:2] != pipe_tx08_eq_control)? 1'b1 : 1'b0; 
  assign pipe_tx09_eq_done = (pipe_tx09_eq_control_reg[3:2] != pipe_tx09_eq_control)? 1'b1 : 1'b0; 
  assign pipe_tx10_eq_done = (pipe_tx10_eq_control_reg[3:2] != pipe_tx10_eq_control)? 1'b1 : 1'b0; 
  assign pipe_tx11_eq_done = (pipe_tx11_eq_control_reg[3:2] != pipe_tx11_eq_control)? 1'b1 : 1'b0; 
  assign pipe_tx12_eq_done = (pipe_tx12_eq_control_reg[3:2] != pipe_tx12_eq_control)? 1'b1 : 1'b0; 
  assign pipe_tx13_eq_done = (pipe_tx13_eq_control_reg[3:2] != pipe_tx13_eq_control)? 1'b1 : 1'b0; 
  assign pipe_tx14_eq_done = (pipe_tx14_eq_control_reg[3:2] != pipe_tx14_eq_control)? 1'b1 : 1'b0; 
  assign pipe_tx15_eq_done = (pipe_tx15_eq_control_reg[3:2] != pipe_tx15_eq_control)? 1'b1 : 1'b0; 
 
 // Pipe mode tie-offs
 assign  common_commands_out[0]    = pipe_clk;
 assign  common_commands_out[3]    = pipe_tx0_rcvr_det; 
 assign  common_commands_out[16:10] = 7'b0;
 assign  pipe_tx_0_sigs[69:42]     = 28'b0;
 assign  pipe_tx_1_sigs[69:42]     = 28'b0;
 assign  pipe_tx_2_sigs[69:42]     = 28'b0;
 assign  pipe_tx_3_sigs[69:42]     = 28'b0;
 assign  pipe_tx_4_sigs[69:42]     = 28'b0;
 assign  pipe_tx_5_sigs[69:42]     = 28'b0;
 assign  pipe_tx_6_sigs[69:42]     = 28'b0;
 assign  pipe_tx_7_sigs[69:42]     = 28'b0; 
 assign  pipe_tx_8_sigs[69:42]     = 28'b0; 
 assign  pipe_tx_9_sigs[69:42]     = 28'b0; 
 assign  pipe_tx_10_sigs[69:42]     = 28'b0; 
 assign  pipe_tx_11_sigs[69:42]     = 28'b0; 
 assign  pipe_tx_12_sigs[69:42]     = 28'b0; 
 assign  pipe_tx_13_sigs[69:42]     = 28'b0; 
 assign  pipe_tx_14_sigs[69:42]     = 28'b0; 
 assign  pipe_tx_15_sigs[69:42]     = 28'b0; 

 end
endgenerate

generate if (EXT_PIPE_SIM == "FALSE") 
begin
  xp4_usp_smsw_pipe 
 #(
    .TCQ(TCQ)
   ,.IMPL_TARGET(IMPL_TARGET)
   ,.AXISTEN_IF_EXT_512_INTFC_RAM_STYLE(AXISTEN_IF_EXT_512_INTFC_RAM_STYLE)
   ,.CRM_CORE_CLK_FREQ_500(CRM_CORE_CLK_FREQ_500)
   ,.CRM_USER_CLK_FREQ(CRM_USER_CLK_FREQ)
   ,.AXISTEN_IF_WIDTH(AXISTEN_IF_WIDTH)
   ,.AXISTEN_IF_EXT_512_CQ_STRADDLE(AXISTEN_IF_EXT_512_CQ_STRADDLE)
   ,.AXISTEN_IF_EXT_512_CC_STRADDLE(AXISTEN_IF_EXT_512_CC_STRADDLE)
   ,.AXISTEN_IF_EXT_512_RQ_STRADDLE(AXISTEN_IF_EXT_512_RQ_STRADDLE)
   ,.AXISTEN_IF_EXT_512_RC_STRADDLE(AXISTEN_IF_EXT_512_RC_STRADDLE)
   ,.AXISTEN_IF_EXT_512_RC_4TLP_STRADDLE(AXISTEN_IF_EXT_512_RC_4TLP_STRADDLE)
   ,.AXISTEN_IF_EXT_512(AXISTEN_IF_EXT_512)
   ,.AXISTEN_IF_CQ_ALIGNMENT_MODE(AXISTEN_IF_CQ_ALIGNMENT_MODE)
   ,.AXISTEN_IF_CC_ALIGNMENT_MODE(AXISTEN_IF_CC_ALIGNMENT_MODE)
   ,.AXISTEN_IF_RQ_ALIGNMENT_MODE(AXISTEN_IF_RQ_ALIGNMENT_MODE)
   ,.AXISTEN_IF_RC_ALIGNMENT_MODE(AXISTEN_IF_RC_ALIGNMENT_MODE)
   ,.AXISTEN_IF_RC_STRADDLE(AXISTEN_IF_RC_STRADDLE)
   ,.AXI4_DATA_WIDTH(AXI4_DATA_WIDTH)
   ,.AXI4_TKEEP_WIDTH(AXI4_TKEEP_WIDTH)
   ,.AXI4_CQ_TUSER_WIDTH(AXI4_CQ_TUSER_WIDTH)
   ,.AXI4_CC_TUSER_WIDTH(AXI4_CC_TUSER_WIDTH)
   ,.AXI4_RQ_TUSER_WIDTH(AXI4_RQ_TUSER_WIDTH)
   ,.AXI4_RC_TUSER_WIDTH(AXI4_RC_TUSER_WIDTH)
   ,.AXI4_CQ_TREADY_WIDTH(AXI4_CQ_TREADY_WIDTH)
   ,.AXI4_CC_TREADY_WIDTH(AXI4_CC_TREADY_WIDTH)
   ,.AXI4_RQ_TREADY_WIDTH(AXI4_RQ_TREADY_WIDTH)
   ,.AXI4_RC_TREADY_WIDTH(AXI4_RC_TREADY_WIDTH)
   ,.AXISTEN_IF_ENABLE_RX_MSG_INTFC(AXISTEN_IF_ENABLE_RX_MSG_INTFC)
   ,.AXISTEN_IF_ENABLE_MSG_ROUTE(AXISTEN_IF_ENABLE_MSG_ROUTE)
   ,.AXISTEN_IF_RX_PARITY_EN(AXISTEN_IF_RX_PARITY_EN)
   ,.AXISTEN_IF_TX_PARITY_EN(AXISTEN_IF_TX_PARITY_EN)
   ,.AXISTEN_IF_ENABLE_CLIENT_TAG(AXISTEN_IF_ENABLE_CLIENT_TAG)
   ,.AXISTEN_IF_ENABLE_256_TAGS(AXISTEN_IF_ENABLE_256_TAGS)
   ,.AXISTEN_IF_COMPL_TIMEOUT_REG0(AXISTEN_IF_COMPL_TIMEOUT_REG0)
   ,.AXISTEN_IF_COMPL_TIMEOUT_REG1(AXISTEN_IF_COMPL_TIMEOUT_REG1)
   ,.AXISTEN_IF_LEGACY_MODE_ENABLE(AXISTEN_IF_LEGACY_MODE_ENABLE)
   ,.AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK(AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK)
   ,.AXISTEN_IF_MSIX_TO_RAM_PIPELINE(AXISTEN_IF_MSIX_TO_RAM_PIPELINE)
   ,.AXISTEN_IF_MSIX_FROM_RAM_PIPELINE(AXISTEN_IF_MSIX_FROM_RAM_PIPELINE)
   ,.AXISTEN_IF_MSIX_RX_PARITY_EN(AXISTEN_IF_MSIX_RX_PARITY_EN)
   ,.AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE(AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE)
   ,.AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT(AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT)
   ,.AXISTEN_IF_CQ_EN_POISONED_MEM_WR(AXISTEN_IF_CQ_EN_POISONED_MEM_WR)
   ,.AXISTEN_IF_RQ_CC_REGISTERED_TREADY(AXISTEN_IF_RQ_CC_REGISTERED_TREADY)
   ,.PM_ASPML0S_TIMEOUT(PM_ASPML0S_TIMEOUT)
   ,.PM_L1_REENTRY_DELAY(PM_L1_REENTRY_DELAY)
   ,.PM_ASPML1_ENTRY_DELAY(PM_ASPML1_ENTRY_DELAY)
   ,.PM_ENABLE_SLOT_POWER_CAPTURE(PM_ENABLE_SLOT_POWER_CAPTURE)
   ,.PM_PME_SERVICE_TIMEOUT_DELAY(PM_PME_SERVICE_TIMEOUT_DELAY)
   ,.PM_PME_TURNOFF_ACK_DELAY(PM_PME_TURNOFF_ACK_DELAY)
   ,.PL_UPSTREAM_FACING(PL_UPSTREAM_FACING)
   ,.PL_LINK_CAP_MAX_LINK_WIDTH(PL_LINK_CAP_MAX_LINK_WIDTH)
   ,.PL_LINK_CAP_MAX_LINK_SPEED(PL_LINK_CAP_MAX_LINK_SPEED)
   ,.PL_DISABLE_DC_BALANCE(PL_DISABLE_DC_BALANCE)
   ,.PL_DISABLE_EI_INFER_IN_L0(PL_DISABLE_EI_INFER_IN_L0)
   ,.PL_N_FTS(PL_N_FTS)
   ,.PL_DISABLE_UPCONFIG_CAPABLE(PL_DISABLE_UPCONFIG_CAPABLE)
   ,.PL_DISABLE_RETRAIN_ON_FRAMING_ERROR(PL_DISABLE_RETRAIN_ON_FRAMING_ERROR)
   ,.PL_DISABLE_RETRAIN_ON_EB_ERROR(PL_DISABLE_RETRAIN_ON_EB_ERROR)
   ,.PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR(PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR)
   ,.PL_REPORT_ALL_PHY_ERRORS(PL_REPORT_ALL_PHY_ERRORS)
   ,.PL_DISABLE_LFSR_UPDATE_ON_SKP(PL_DISABLE_LFSR_UPDATE_ON_SKP)
   ,.PL_LANE0_EQ_CONTROL(PL_LANE0_EQ_CONTROL)
   ,.PL_LANE1_EQ_CONTROL(PL_LANE1_EQ_CONTROL)
   ,.PL_LANE2_EQ_CONTROL(PL_LANE2_EQ_CONTROL)
   ,.PL_LANE3_EQ_CONTROL(PL_LANE3_EQ_CONTROL)
   ,.PL_LANE4_EQ_CONTROL(PL_LANE4_EQ_CONTROL)
   ,.PL_LANE5_EQ_CONTROL(PL_LANE5_EQ_CONTROL)
   ,.PL_LANE6_EQ_CONTROL(PL_LANE6_EQ_CONTROL)
   ,.PL_LANE7_EQ_CONTROL(PL_LANE7_EQ_CONTROL)
   ,.PL_LANE8_EQ_CONTROL(PL_LANE8_EQ_CONTROL)
   ,.PL_LANE9_EQ_CONTROL(PL_LANE9_EQ_CONTROL)
   ,.PL_LANE10_EQ_CONTROL(PL_LANE10_EQ_CONTROL)
   ,.PL_LANE11_EQ_CONTROL(PL_LANE11_EQ_CONTROL)
   ,.PL_LANE12_EQ_CONTROL(PL_LANE12_EQ_CONTROL)
   ,.PL_LANE13_EQ_CONTROL(PL_LANE13_EQ_CONTROL)
   ,.PL_LANE14_EQ_CONTROL(PL_LANE14_EQ_CONTROL)
   ,.PL_LANE15_EQ_CONTROL(PL_LANE15_EQ_CONTROL)
   ,.PL_EQ_BYPASS_PHASE23(PL_EQ_BYPASS_PHASE23)
   ,.PL_EQ_ADAPT_ITER_COUNT(PL_EQ_ADAPT_ITER_COUNT)
   ,.PL_EQ_ADAPT_REJECT_RETRY_COUNT(PL_EQ_ADAPT_REJECT_RETRY_COUNT)
   ,.PL_EQ_SHORT_ADAPT_PHASE(PL_EQ_SHORT_ADAPT_PHASE)
   ,.PL_EQ_ADAPT_DISABLE_COEFF_CHECK(PL_EQ_ADAPT_DISABLE_COEFF_CHECK)
   ,.PL_EQ_ADAPT_DISABLE_PRESET_CHECK(PL_EQ_ADAPT_DISABLE_PRESET_CHECK)
   ,.PL_EQ_DEFAULT_TX_PRESET(PL_EQ_DEFAULT_TX_PRESET)
   ,.PL_EQ_DEFAULT_RX_PRESET_HINT(PL_EQ_DEFAULT_RX_PRESET_HINT)
   ,.PL_EQ_RX_ADAPT_EQ_PHASE0(PL_EQ_RX_ADAPT_EQ_PHASE0)
   ,.PL_EQ_RX_ADAPT_EQ_PHASE1(PL_EQ_RX_ADAPT_EQ_PHASE1)
   ,.PL_EQ_DISABLE_MISMATCH_CHECK(PL_EQ_DISABLE_MISMATCH_CHECK)
   ,.PL_RX_L0S_EXIT_TO_RECOVERY(PL_RX_L0S_EXIT_TO_RECOVERY)
   ,.PL_EQ_TX_8G_EQ_TS2_ENABLE(PL_EQ_TX_8G_EQ_TS2_ENABLE)
   ,.PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4(PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4)
   ,.PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3(PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3)
   ,.PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2(PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2)
   ,.PL_DESKEW_ON_SKIP_IN_GEN12(PL_DESKEW_ON_SKIP_IN_GEN12)
   ,.PL_INFER_EI_DISABLE_REC_RC(PL_INFER_EI_DISABLE_REC_RC)
   ,.PL_INFER_EI_DISABLE_REC_SPD(PL_INFER_EI_DISABLE_REC_SPD)
   ,.PL_INFER_EI_DISABLE_LPBK_ACTIVE(PL_INFER_EI_DISABLE_LPBK_ACTIVE)
   ,.PL_RX_ADAPT_TIMER_RRL_GEN3(PL_RX_ADAPT_TIMER_RRL_GEN3)
   ,.PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS(PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS)
   ,.PL_RX_ADAPT_TIMER_RRL_GEN4(PL_RX_ADAPT_TIMER_RRL_GEN4)
   ,.PL_RX_ADAPT_TIMER_CLWS_GEN3(PL_RX_ADAPT_TIMER_CLWS_GEN3)
   ,.PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS(PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS)
   ,.PL_RX_ADAPT_TIMER_CLWS_GEN4(PL_RX_ADAPT_TIMER_CLWS_GEN4)
   ,.PL_DISABLE_LANE_REVERSAL(PL_DISABLE_LANE_REVERSAL)
   ,.PL_CFG_STATE_ROBUSTNESS_ENABLE(PL_CFG_STATE_ROBUSTNESS_ENABLE)
   ,.PL_REDO_EQ_SOURCE_SELECT(PL_REDO_EQ_SOURCE_SELECT)
   ,.PL_DEEMPH_SOURCE_SELECT(PL_DEEMPH_SOURCE_SELECT)
   ,.PL_EXIT_LOOPBACK_ON_EI_ENTRY(PL_EXIT_LOOPBACK_ON_EI_ENTRY)
   ,.PL_QUIESCE_GUARANTEE_DISABLE(PL_QUIESCE_GUARANTEE_DISABLE)
   ,.PL_SRIS_ENABLE(PL_SRIS_ENABLE)
   ,.PL_SRIS_SKPOS_GEN_SPD_VEC(PL_SRIS_SKPOS_GEN_SPD_VEC)
   ,.PL_SRIS_SKPOS_REC_SPD_VEC(PL_SRIS_SKPOS_REC_SPD_VEC)
   ,.PL_SIM_FAST_LINK_TRAINING(PL_SIM_FAST_LINK_TRAINING)
   ,.PL_USER_SPARE(PL_USER_SPARE)
   ,.LL_ACK_TIMEOUT_EN(LL_ACK_TIMEOUT_EN)
   ,.LL_ACK_TIMEOUT(LL_ACK_TIMEOUT)
   ,.LL_ACK_TIMEOUT_FUNC(LL_ACK_TIMEOUT_FUNC)
   ,.LL_REPLAY_TIMEOUT_EN(LL_REPLAY_TIMEOUT_EN)
   ,.LL_REPLAY_TIMEOUT(LL_REPLAY_TIMEOUT)
   ,.LL_REPLAY_TIMEOUT_FUNC(LL_REPLAY_TIMEOUT_FUNC)
   ,.LL_REPLAY_TO_RAM_PIPELINE(LL_REPLAY_TO_RAM_PIPELINE)
   ,.LL_REPLAY_FROM_RAM_PIPELINE(LL_REPLAY_FROM_RAM_PIPELINE)
   ,.LL_DISABLE_SCHED_TX_NAK(LL_DISABLE_SCHED_TX_NAK)
   ,.LL_TX_TLP_PARITY_CHK(LL_TX_TLP_PARITY_CHK)
   ,.LL_RX_TLP_PARITY_GEN(LL_RX_TLP_PARITY_GEN)
   ,.LL_USER_SPARE(LL_USER_SPARE)
   ,.IS_SWITCH_PORT(IS_SWITCH_PORT)
   ,.CFG_BYPASS_MODE_ENABLE(CFG_BYPASS_MODE_ENABLE)
   ,.TL_PF_ENABLE_REG(TL_PF_ENABLE_REG)
   ,.TL_CREDITS_CD(TL_CREDITS_CD)
   ,.TL_CREDITS_CH(TL_CREDITS_CH)
   ,.TL_COMPLETION_RAM_SIZE(TL_COMPLETION_RAM_SIZE)
   ,.TL_COMPLETION_RAM_NUM_TLPS(TL_COMPLETION_RAM_NUM_TLPS)
   ,.TL_CREDITS_NPD(TL_CREDITS_NPD)
   ,.TL_CREDITS_NPH(TL_CREDITS_NPH)
   ,.TL_CREDITS_PD(TL_CREDITS_PD)
   ,.TL_CREDITS_PH(TL_CREDITS_PH)
   ,.TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE(TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE)
   ,.TL_RX_COMPLETION_TO_RAM_READ_PIPELINE(TL_RX_COMPLETION_TO_RAM_READ_PIPELINE)
   ,.TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE(TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE)
   ,.TL_POSTED_RAM_SIZE(TL_POSTED_RAM_SIZE)
   ,.TL_RX_POSTED_TO_RAM_WRITE_PIPELINE(TL_RX_POSTED_TO_RAM_WRITE_PIPELINE)
   ,.TL_RX_POSTED_TO_RAM_READ_PIPELINE(TL_RX_POSTED_TO_RAM_READ_PIPELINE)
   ,.TL_RX_POSTED_FROM_RAM_READ_PIPELINE(TL_RX_POSTED_FROM_RAM_READ_PIPELINE)
   ,.TL_TX_MUX_STRICT_PRIORITY(TL_TX_MUX_STRICT_PRIORITY)
   ,.TL_TX_TLP_STRADDLE_ENABLE(TL_TX_TLP_STRADDLE_ENABLE)
   ,.TL_TX_TLP_TERMINATE_PARITY(TL_TX_TLP_TERMINATE_PARITY)
   ,.TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT(TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT)
   ,.TL_FC_UPDATE_MIN_INTERVAL_TIME(TL_FC_UPDATE_MIN_INTERVAL_TIME)
   ,.TL_USER_SPARE(TL_USER_SPARE)
   ,.PF0_CLASS_CODE(PF0_CLASS_CODE)
   ,.PF1_CLASS_CODE(PF1_CLASS_CODE)
   ,.PF2_CLASS_CODE(PF2_CLASS_CODE)
   ,.PF3_CLASS_CODE(PF3_CLASS_CODE)
   ,.PF0_INTERRUPT_PIN(PF0_INTERRUPT_PIN)
   ,.PF1_INTERRUPT_PIN(PF1_INTERRUPT_PIN)
   ,.PF2_INTERRUPT_PIN(PF2_INTERRUPT_PIN)
   ,.PF3_INTERRUPT_PIN(PF3_INTERRUPT_PIN)
   ,.PF0_CAPABILITY_POINTER(PF0_CAPABILITY_POINTER)
   ,.PF1_CAPABILITY_POINTER(PF1_CAPABILITY_POINTER)
   ,.PF2_CAPABILITY_POINTER(PF2_CAPABILITY_POINTER)
   ,.PF3_CAPABILITY_POINTER(PF3_CAPABILITY_POINTER)
   ,.VF0_CAPABILITY_POINTER(VF0_CAPABILITY_POINTER)
   ,.LEGACY_CFG_EXTEND_INTERFACE_ENABLE(LEGACY_CFG_EXTEND_INTERFACE_ENABLE)
   ,.EXTENDED_CFG_EXTEND_INTERFACE_ENABLE(EXTENDED_CFG_EXTEND_INTERFACE_ENABLE)
   ,.TL2CFG_IF_PARITY_CHK(TL2CFG_IF_PARITY_CHK)
   ,.HEADER_TYPE_OVERRIDE(HEADER_TYPE_OVERRIDE)
   ,.PF0_BAR0_CONTROL(PF0_BAR0_CONTROL)
   ,.PF1_BAR0_CONTROL(PF1_BAR0_CONTROL)
   ,.PF2_BAR0_CONTROL(PF2_BAR0_CONTROL)
   ,.PF3_BAR0_CONTROL(PF3_BAR0_CONTROL)
   ,.PF0_BAR0_APERTURE_SIZE(PF0_BAR0_APERTURE_SIZE)
   ,.PF1_BAR0_APERTURE_SIZE(PF1_BAR0_APERTURE_SIZE)
   ,.PF2_BAR0_APERTURE_SIZE(PF2_BAR0_APERTURE_SIZE)
   ,.PF3_BAR0_APERTURE_SIZE(PF3_BAR0_APERTURE_SIZE)
   ,.PF0_BAR1_CONTROL(PF0_BAR1_CONTROL)
   ,.PF1_BAR1_CONTROL(PF1_BAR1_CONTROL)
   ,.PF2_BAR1_CONTROL(PF2_BAR1_CONTROL)
   ,.PF3_BAR1_CONTROL(PF3_BAR1_CONTROL)
   ,.PF0_BAR1_APERTURE_SIZE(PF0_BAR1_APERTURE_SIZE)
   ,.PF1_BAR1_APERTURE_SIZE(PF1_BAR1_APERTURE_SIZE)
   ,.PF2_BAR1_APERTURE_SIZE(PF2_BAR1_APERTURE_SIZE)
   ,.PF3_BAR1_APERTURE_SIZE(PF3_BAR1_APERTURE_SIZE)
   ,.PF0_BAR2_CONTROL(PF0_BAR2_CONTROL)
   ,.PF1_BAR2_CONTROL(PF1_BAR2_CONTROL)
   ,.PF2_BAR2_CONTROL(PF2_BAR2_CONTROL)
   ,.PF3_BAR2_CONTROL(PF3_BAR2_CONTROL)
   ,.PF0_BAR2_APERTURE_SIZE(PF0_BAR2_APERTURE_SIZE)
   ,.PF1_BAR2_APERTURE_SIZE(PF1_BAR2_APERTURE_SIZE)
   ,.PF2_BAR2_APERTURE_SIZE(PF2_BAR2_APERTURE_SIZE)
   ,.PF3_BAR2_APERTURE_SIZE(PF3_BAR2_APERTURE_SIZE)
   ,.PF0_BAR3_CONTROL(PF0_BAR3_CONTROL)
   ,.PF1_BAR3_CONTROL(PF1_BAR3_CONTROL)
   ,.PF2_BAR3_CONTROL(PF2_BAR3_CONTROL)
   ,.PF3_BAR3_CONTROL(PF3_BAR3_CONTROL)
   ,.PF0_BAR3_APERTURE_SIZE(PF0_BAR3_APERTURE_SIZE)
   ,.PF1_BAR3_APERTURE_SIZE(PF1_BAR3_APERTURE_SIZE)
   ,.PF2_BAR3_APERTURE_SIZE(PF2_BAR3_APERTURE_SIZE)
   ,.PF3_BAR3_APERTURE_SIZE(PF3_BAR3_APERTURE_SIZE)
   ,.PF0_BAR4_CONTROL(PF0_BAR4_CONTROL)
   ,.PF1_BAR4_CONTROL(PF1_BAR4_CONTROL)
   ,.PF2_BAR4_CONTROL(PF2_BAR4_CONTROL)
   ,.PF3_BAR4_CONTROL(PF3_BAR4_CONTROL)
   ,.PF0_BAR4_APERTURE_SIZE(PF0_BAR4_APERTURE_SIZE)
   ,.PF1_BAR4_APERTURE_SIZE(PF1_BAR4_APERTURE_SIZE)
   ,.PF2_BAR4_APERTURE_SIZE(PF2_BAR4_APERTURE_SIZE)
   ,.PF3_BAR4_APERTURE_SIZE(PF3_BAR4_APERTURE_SIZE)
   ,.PF0_BAR5_CONTROL(PF0_BAR5_CONTROL)
   ,.PF1_BAR5_CONTROL(PF1_BAR5_CONTROL)
   ,.PF2_BAR5_CONTROL(PF2_BAR5_CONTROL)
   ,.PF3_BAR5_CONTROL(PF3_BAR5_CONTROL)
   ,.PF0_BAR5_APERTURE_SIZE(PF0_BAR5_APERTURE_SIZE)
   ,.PF1_BAR5_APERTURE_SIZE(PF1_BAR5_APERTURE_SIZE)
   ,.PF2_BAR5_APERTURE_SIZE(PF2_BAR5_APERTURE_SIZE)
   ,.PF3_BAR5_APERTURE_SIZE(PF3_BAR5_APERTURE_SIZE)
   ,.PF0_EXPANSION_ROM_ENABLE(PF0_EXPANSION_ROM_ENABLE)
   ,.PF1_EXPANSION_ROM_ENABLE(PF1_EXPANSION_ROM_ENABLE)
   ,.PF2_EXPANSION_ROM_ENABLE(PF2_EXPANSION_ROM_ENABLE)
   ,.PF3_EXPANSION_ROM_ENABLE(PF3_EXPANSION_ROM_ENABLE)
   ,.PF0_EXPANSION_ROM_APERTURE_SIZE(PF0_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF1_EXPANSION_ROM_APERTURE_SIZE(PF1_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF2_EXPANSION_ROM_APERTURE_SIZE(PF2_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF3_EXPANSION_ROM_APERTURE_SIZE(PF3_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF0_PCIE_CAP_NEXTPTR(PF0_PCIE_CAP_NEXTPTR)
   ,.PF1_PCIE_CAP_NEXTPTR(PF1_PCIE_CAP_NEXTPTR)
   ,.PF2_PCIE_CAP_NEXTPTR(PF2_PCIE_CAP_NEXTPTR)
   ,.PF3_PCIE_CAP_NEXTPTR(PF3_PCIE_CAP_NEXTPTR)
   ,.VFG0_PCIE_CAP_NEXTPTR(VFG0_PCIE_CAP_NEXTPTR)
   ,.VFG1_PCIE_CAP_NEXTPTR(VFG1_PCIE_CAP_NEXTPTR)
   ,.VFG2_PCIE_CAP_NEXTPTR(VFG2_PCIE_CAP_NEXTPTR)
   ,.VFG3_PCIE_CAP_NEXTPTR(VFG3_PCIE_CAP_NEXTPTR)
   ,.PF0_DEV_CAP_MAX_PAYLOAD_SIZE(PF0_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF1_DEV_CAP_MAX_PAYLOAD_SIZE(PF1_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF2_DEV_CAP_MAX_PAYLOAD_SIZE(PF2_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF3_DEV_CAP_MAX_PAYLOAD_SIZE(PF3_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF0_DEV_CAP_EXT_TAG_SUPPORTED(PF0_DEV_CAP_EXT_TAG_SUPPORTED)
   ,.PF0_DEV_CAP_ENDPOINT_L0S_LATENCY(PF0_DEV_CAP_ENDPOINT_L0S_LATENCY)
   ,.PF0_DEV_CAP_ENDPOINT_L1_LATENCY(PF0_DEV_CAP_ENDPOINT_L1_LATENCY)
   ,.PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE(PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE)
   ,.PF0_LINK_CAP_ASPM_SUPPORT(PF0_LINK_CAP_ASPM_SUPPORT)
   ,.PF0_LINK_CONTROL_RCB(PF0_LINK_CONTROL_RCB)
   ,.PF0_LINK_STATUS_SLOT_CLOCK_CONFIG(PF0_LINK_STATUS_SLOT_CLOCK_CONFIG)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4)
   ,.PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE(PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE)
   ,.PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT(PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT(PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT(PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_LTR_SUPPORT(PF0_DEV_CAP2_LTR_SUPPORT)
   ,.PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT(PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_OBFF_SUPPORT(PF0_DEV_CAP2_OBFF_SUPPORT)
   ,.PF0_DEV_CAP2_ARI_FORWARD_ENABLE(PF0_DEV_CAP2_ARI_FORWARD_ENABLE)
   ,.PF0_MSI_CAP_NEXTPTR(PF0_MSI_CAP_NEXTPTR)
   ,.PF1_MSI_CAP_NEXTPTR(PF1_MSI_CAP_NEXTPTR)
   ,.PF2_MSI_CAP_NEXTPTR(PF2_MSI_CAP_NEXTPTR)
   ,.PF3_MSI_CAP_NEXTPTR(PF3_MSI_CAP_NEXTPTR)
   ,.PF0_MSI_CAP_PERVECMASKCAP(PF0_MSI_CAP_PERVECMASKCAP)
   ,.PF1_MSI_CAP_PERVECMASKCAP(PF1_MSI_CAP_PERVECMASKCAP)
   ,.PF2_MSI_CAP_PERVECMASKCAP(PF2_MSI_CAP_PERVECMASKCAP)
   ,.PF3_MSI_CAP_PERVECMASKCAP(PF3_MSI_CAP_PERVECMASKCAP)
   ,.PF0_MSI_CAP_MULTIMSGCAP(PF0_MSI_CAP_MULTIMSGCAP)
   ,.PF1_MSI_CAP_MULTIMSGCAP(PF1_MSI_CAP_MULTIMSGCAP)
   ,.PF2_MSI_CAP_MULTIMSGCAP(PF2_MSI_CAP_MULTIMSGCAP)
   ,.PF3_MSI_CAP_MULTIMSGCAP(PF3_MSI_CAP_MULTIMSGCAP)
   ,.PF0_MSIX_CAP_NEXTPTR(PF0_MSIX_CAP_NEXTPTR)
   ,.PF1_MSIX_CAP_NEXTPTR(PF1_MSIX_CAP_NEXTPTR)
   ,.PF2_MSIX_CAP_NEXTPTR(PF2_MSIX_CAP_NEXTPTR)
   ,.PF3_MSIX_CAP_NEXTPTR(PF3_MSIX_CAP_NEXTPTR)
   ,.VFG0_MSIX_CAP_NEXTPTR(VFG0_MSIX_CAP_NEXTPTR)
   ,.VFG1_MSIX_CAP_NEXTPTR(VFG1_MSIX_CAP_NEXTPTR)
   ,.VFG2_MSIX_CAP_NEXTPTR(VFG2_MSIX_CAP_NEXTPTR)
   ,.VFG3_MSIX_CAP_NEXTPTR(VFG3_MSIX_CAP_NEXTPTR)
   ,.PF0_MSIX_CAP_PBA_BIR(PF0_MSIX_CAP_PBA_BIR)
   ,.PF1_MSIX_CAP_PBA_BIR(PF1_MSIX_CAP_PBA_BIR)
   ,.PF2_MSIX_CAP_PBA_BIR(PF2_MSIX_CAP_PBA_BIR)
   ,.PF3_MSIX_CAP_PBA_BIR(PF3_MSIX_CAP_PBA_BIR)
   ,.VFG0_MSIX_CAP_PBA_BIR(VFG0_MSIX_CAP_PBA_BIR)
   ,.VFG1_MSIX_CAP_PBA_BIR(VFG1_MSIX_CAP_PBA_BIR)
   ,.VFG2_MSIX_CAP_PBA_BIR(VFG2_MSIX_CAP_PBA_BIR)
   ,.VFG3_MSIX_CAP_PBA_BIR(VFG3_MSIX_CAP_PBA_BIR)
   ,.PF0_MSIX_CAP_PBA_OFFSET(PF0_MSIX_CAP_PBA_OFFSET)
   ,.PF1_MSIX_CAP_PBA_OFFSET(PF1_MSIX_CAP_PBA_OFFSET)
   ,.PF2_MSIX_CAP_PBA_OFFSET(PF2_MSIX_CAP_PBA_OFFSET)
   ,.PF3_MSIX_CAP_PBA_OFFSET(PF3_MSIX_CAP_PBA_OFFSET)
   ,.VFG0_MSIX_CAP_PBA_OFFSET(VFG0_MSIX_CAP_PBA_OFFSET)
   ,.VFG1_MSIX_CAP_PBA_OFFSET(VFG1_MSIX_CAP_PBA_OFFSET)
   ,.VFG2_MSIX_CAP_PBA_OFFSET(VFG2_MSIX_CAP_PBA_OFFSET)
   ,.VFG3_MSIX_CAP_PBA_OFFSET(VFG3_MSIX_CAP_PBA_OFFSET)
   ,.PF0_MSIX_CAP_TABLE_BIR(PF0_MSIX_CAP_TABLE_BIR)
   ,.PF1_MSIX_CAP_TABLE_BIR(PF1_MSIX_CAP_TABLE_BIR)
   ,.PF2_MSIX_CAP_TABLE_BIR(PF2_MSIX_CAP_TABLE_BIR)
   ,.PF3_MSIX_CAP_TABLE_BIR(PF3_MSIX_CAP_TABLE_BIR)
   ,.VFG0_MSIX_CAP_TABLE_BIR(VFG0_MSIX_CAP_TABLE_BIR)
   ,.VFG1_MSIX_CAP_TABLE_BIR(VFG1_MSIX_CAP_TABLE_BIR)
   ,.VFG2_MSIX_CAP_TABLE_BIR(VFG2_MSIX_CAP_TABLE_BIR)
   ,.VFG3_MSIX_CAP_TABLE_BIR(VFG3_MSIX_CAP_TABLE_BIR)
   ,.PF0_MSIX_CAP_TABLE_OFFSET(PF0_MSIX_CAP_TABLE_OFFSET)
   ,.PF1_MSIX_CAP_TABLE_OFFSET(PF1_MSIX_CAP_TABLE_OFFSET)
   ,.PF2_MSIX_CAP_TABLE_OFFSET(PF2_MSIX_CAP_TABLE_OFFSET)
   ,.PF3_MSIX_CAP_TABLE_OFFSET(PF3_MSIX_CAP_TABLE_OFFSET)
   ,.VFG0_MSIX_CAP_TABLE_OFFSET(VFG0_MSIX_CAP_TABLE_OFFSET)
   ,.VFG1_MSIX_CAP_TABLE_OFFSET(VFG1_MSIX_CAP_TABLE_OFFSET)
   ,.VFG2_MSIX_CAP_TABLE_OFFSET(VFG2_MSIX_CAP_TABLE_OFFSET)
   ,.VFG3_MSIX_CAP_TABLE_OFFSET(VFG3_MSIX_CAP_TABLE_OFFSET)
   ,.PF0_MSIX_CAP_TABLE_SIZE(PF0_MSIX_CAP_TABLE_SIZE)
   ,.PF1_MSIX_CAP_TABLE_SIZE(PF1_MSIX_CAP_TABLE_SIZE)
   ,.PF2_MSIX_CAP_TABLE_SIZE(PF2_MSIX_CAP_TABLE_SIZE)
   ,.PF3_MSIX_CAP_TABLE_SIZE(PF3_MSIX_CAP_TABLE_SIZE)
   ,.VFG0_MSIX_CAP_TABLE_SIZE(VFG0_MSIX_CAP_TABLE_SIZE)
   ,.VFG1_MSIX_CAP_TABLE_SIZE(VFG1_MSIX_CAP_TABLE_SIZE)
   ,.VFG2_MSIX_CAP_TABLE_SIZE(VFG2_MSIX_CAP_TABLE_SIZE)
   ,.VFG3_MSIX_CAP_TABLE_SIZE(VFG3_MSIX_CAP_TABLE_SIZE)
   ,.PF0_MSIX_VECTOR_COUNT(PF0_MSIX_VECTOR_COUNT)
   ,.PF0_PM_CAP_ID(PF0_PM_CAP_ID)
   ,.PF0_PM_CAP_NEXTPTR(PF0_PM_CAP_NEXTPTR)
   ,.PF1_PM_CAP_NEXTPTR(PF1_PM_CAP_NEXTPTR)
   ,.PF2_PM_CAP_NEXTPTR(PF2_PM_CAP_NEXTPTR)
   ,.PF3_PM_CAP_NEXTPTR(PF3_PM_CAP_NEXTPTR)
   ,.PF0_PM_CAP_PMESUPPORT_D3HOT(PF0_PM_CAP_PMESUPPORT_D3HOT)
   ,.PF0_PM_CAP_PMESUPPORT_D1(PF0_PM_CAP_PMESUPPORT_D1)
   ,.PF0_PM_CAP_PMESUPPORT_D0(PF0_PM_CAP_PMESUPPORT_D0)
   ,.PF0_PM_CAP_SUPP_D1_STATE(PF0_PM_CAP_SUPP_D1_STATE)
   ,.PF0_PM_CAP_VER_ID(PF0_PM_CAP_VER_ID)
   ,.PF0_PM_CSR_NOSOFTRESET(PF0_PM_CSR_NOSOFTRESET)
   ,.PM_ENABLE_L23_ENTRY(PM_ENABLE_L23_ENTRY)
   ,.DNSTREAM_LINK_NUM(DNSTREAM_LINK_NUM)
   ,.AUTO_FLR_RESPONSE(AUTO_FLR_RESPONSE)
   ,.PF0_DSN_CAP_NEXTPTR(PF0_DSN_CAP_NEXTPTR)
   ,.PF1_DSN_CAP_NEXTPTR(PF1_DSN_CAP_NEXTPTR)
   ,.PF2_DSN_CAP_NEXTPTR(PF2_DSN_CAP_NEXTPTR)
   ,.PF3_DSN_CAP_NEXTPTR(PF3_DSN_CAP_NEXTPTR)
   ,.DSN_CAP_ENABLE(DSN_CAP_ENABLE)
   ,.PF0_VC_CAP_VER(PF0_VC_CAP_VER)
   ,.PF0_VC_CAP_NEXTPTR(PF0_VC_CAP_NEXTPTR)
   ,.PF0_VC_CAP_ENABLE(PF0_VC_CAP_ENABLE)
   ,.PF0_SECONDARY_PCIE_CAP_NEXTPTR(PF0_SECONDARY_PCIE_CAP_NEXTPTR)
   ,.PF0_AER_CAP_NEXTPTR(PF0_AER_CAP_NEXTPTR)
   ,.PF1_AER_CAP_NEXTPTR(PF1_AER_CAP_NEXTPTR)
   ,.PF2_AER_CAP_NEXTPTR(PF2_AER_CAP_NEXTPTR)
   ,.PF3_AER_CAP_NEXTPTR(PF3_AER_CAP_NEXTPTR)
   ,.PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE(PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE)
   ,.ARI_CAP_ENABLE(ARI_CAP_ENABLE)
   ,.PF0_ARI_CAP_NEXTPTR(PF0_ARI_CAP_NEXTPTR)
   ,.PF1_ARI_CAP_NEXTPTR(PF1_ARI_CAP_NEXTPTR)
   ,.PF2_ARI_CAP_NEXTPTR(PF2_ARI_CAP_NEXTPTR)
   ,.PF3_ARI_CAP_NEXTPTR(PF3_ARI_CAP_NEXTPTR)
   ,.VFG0_ARI_CAP_NEXTPTR(VFG0_ARI_CAP_NEXTPTR)
   ,.VFG1_ARI_CAP_NEXTPTR(VFG1_ARI_CAP_NEXTPTR)
   ,.VFG2_ARI_CAP_NEXTPTR(VFG2_ARI_CAP_NEXTPTR)
   ,.VFG3_ARI_CAP_NEXTPTR(VFG3_ARI_CAP_NEXTPTR)
   ,.PF0_ARI_CAP_VER(PF0_ARI_CAP_VER)
   ,.PF0_ARI_CAP_NEXT_FUNC(PF0_ARI_CAP_NEXT_FUNC)
   ,.PF1_ARI_CAP_NEXT_FUNC(PF1_ARI_CAP_NEXT_FUNC)
   ,.PF2_ARI_CAP_NEXT_FUNC(PF2_ARI_CAP_NEXT_FUNC)
   ,.PF3_ARI_CAP_NEXT_FUNC(PF3_ARI_CAP_NEXT_FUNC)
   ,.PF0_LTR_CAP_NEXTPTR(PF0_LTR_CAP_NEXTPTR)
   ,.PF0_LTR_CAP_VER(PF0_LTR_CAP_VER)
   ,.PF0_LTR_CAP_MAX_SNOOP_LAT(PF0_LTR_CAP_MAX_SNOOP_LAT)
   ,.PF0_LTR_CAP_MAX_NOSNOOP_LAT(PF0_LTR_CAP_MAX_NOSNOOP_LAT)
   ,.LTR_TX_MESSAGE_ON_LTR_ENABLE(LTR_TX_MESSAGE_ON_LTR_ENABLE)
   ,.LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE(LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE)
   ,.LTR_TX_MESSAGE_MINIMUM_INTERVAL(LTR_TX_MESSAGE_MINIMUM_INTERVAL)
   ,.SRIOV_CAP_ENABLE(SRIOV_CAP_ENABLE)
   ,.PF0_SRIOV_CAP_NEXTPTR(PF0_SRIOV_CAP_NEXTPTR)
   ,.PF1_SRIOV_CAP_NEXTPTR(PF1_SRIOV_CAP_NEXTPTR)
   ,.PF2_SRIOV_CAP_NEXTPTR(PF2_SRIOV_CAP_NEXTPTR)
   ,.PF3_SRIOV_CAP_NEXTPTR(PF3_SRIOV_CAP_NEXTPTR)
   ,.PF0_SRIOV_CAP_VER(PF0_SRIOV_CAP_VER)
   ,.PF1_SRIOV_CAP_VER(PF1_SRIOV_CAP_VER)
   ,.PF2_SRIOV_CAP_VER(PF2_SRIOV_CAP_VER)
   ,.PF3_SRIOV_CAP_VER(PF3_SRIOV_CAP_VER)
   ,.PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF0_SRIOV_CAP_INITIAL_VF(PF0_SRIOV_CAP_INITIAL_VF)
   ,.PF1_SRIOV_CAP_INITIAL_VF(PF1_SRIOV_CAP_INITIAL_VF)
   ,.PF2_SRIOV_CAP_INITIAL_VF(PF2_SRIOV_CAP_INITIAL_VF)
   ,.PF3_SRIOV_CAP_INITIAL_VF(PF3_SRIOV_CAP_INITIAL_VF)
   ,.PF0_SRIOV_CAP_TOTAL_VF(PF0_SRIOV_CAP_TOTAL_VF)
   ,.PF1_SRIOV_CAP_TOTAL_VF(PF1_SRIOV_CAP_TOTAL_VF)
   ,.PF2_SRIOV_CAP_TOTAL_VF(PF2_SRIOV_CAP_TOTAL_VF)
   ,.PF3_SRIOV_CAP_TOTAL_VF(PF3_SRIOV_CAP_TOTAL_VF)
   ,.PF0_SRIOV_FUNC_DEP_LINK(PF0_SRIOV_FUNC_DEP_LINK)
   ,.PF1_SRIOV_FUNC_DEP_LINK(PF1_SRIOV_FUNC_DEP_LINK)
   ,.PF2_SRIOV_FUNC_DEP_LINK(PF2_SRIOV_FUNC_DEP_LINK)
   ,.PF3_SRIOV_FUNC_DEP_LINK(PF3_SRIOV_FUNC_DEP_LINK)
   ,.PF0_SRIOV_FIRST_VF_OFFSET(PF0_SRIOV_FIRST_VF_OFFSET)
   ,.PF1_SRIOV_FIRST_VF_OFFSET(PF1_SRIOV_FIRST_VF_OFFSET)
   ,.PF2_SRIOV_FIRST_VF_OFFSET(PF2_SRIOV_FIRST_VF_OFFSET)
   ,.PF3_SRIOV_FIRST_VF_OFFSET(PF3_SRIOV_FIRST_VF_OFFSET)
   ,.PF0_SRIOV_VF_DEVICE_ID(PF0_SRIOV_VF_DEVICE_ID)
   ,.PF1_SRIOV_VF_DEVICE_ID(PF1_SRIOV_VF_DEVICE_ID)
   ,.PF2_SRIOV_VF_DEVICE_ID(PF2_SRIOV_VF_DEVICE_ID)
   ,.PF3_SRIOV_VF_DEVICE_ID(PF3_SRIOV_VF_DEVICE_ID)
   ,.PF0_SRIOV_SUPPORTED_PAGE_SIZE(PF0_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF1_SRIOV_SUPPORTED_PAGE_SIZE(PF1_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF2_SRIOV_SUPPORTED_PAGE_SIZE(PF2_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF3_SRIOV_SUPPORTED_PAGE_SIZE(PF3_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF0_SRIOV_BAR0_CONTROL(PF0_SRIOV_BAR0_CONTROL)
   ,.PF1_SRIOV_BAR0_CONTROL(PF1_SRIOV_BAR0_CONTROL)
   ,.PF2_SRIOV_BAR0_CONTROL(PF2_SRIOV_BAR0_CONTROL)
   ,.PF3_SRIOV_BAR0_CONTROL(PF3_SRIOV_BAR0_CONTROL)
   ,.PF0_SRIOV_BAR0_APERTURE_SIZE(PF0_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR0_APERTURE_SIZE(PF1_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR0_APERTURE_SIZE(PF2_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR0_APERTURE_SIZE(PF3_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR1_CONTROL(PF0_SRIOV_BAR1_CONTROL)
   ,.PF1_SRIOV_BAR1_CONTROL(PF1_SRIOV_BAR1_CONTROL)
   ,.PF2_SRIOV_BAR1_CONTROL(PF2_SRIOV_BAR1_CONTROL)
   ,.PF3_SRIOV_BAR1_CONTROL(PF3_SRIOV_BAR1_CONTROL)
   ,.PF0_SRIOV_BAR1_APERTURE_SIZE(PF0_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR1_APERTURE_SIZE(PF1_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR1_APERTURE_SIZE(PF2_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR1_APERTURE_SIZE(PF3_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR2_CONTROL(PF0_SRIOV_BAR2_CONTROL)
   ,.PF1_SRIOV_BAR2_CONTROL(PF1_SRIOV_BAR2_CONTROL)
   ,.PF2_SRIOV_BAR2_CONTROL(PF2_SRIOV_BAR2_CONTROL)
   ,.PF3_SRIOV_BAR2_CONTROL(PF3_SRIOV_BAR2_CONTROL)
   ,.PF0_SRIOV_BAR2_APERTURE_SIZE(PF0_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR2_APERTURE_SIZE(PF1_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR2_APERTURE_SIZE(PF2_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR2_APERTURE_SIZE(PF3_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR3_CONTROL(PF0_SRIOV_BAR3_CONTROL)
   ,.PF1_SRIOV_BAR3_CONTROL(PF1_SRIOV_BAR3_CONTROL)
   ,.PF2_SRIOV_BAR3_CONTROL(PF2_SRIOV_BAR3_CONTROL)
   ,.PF3_SRIOV_BAR3_CONTROL(PF3_SRIOV_BAR3_CONTROL)
   ,.PF0_SRIOV_BAR3_APERTURE_SIZE(PF0_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR3_APERTURE_SIZE(PF1_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR3_APERTURE_SIZE(PF2_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR3_APERTURE_SIZE(PF3_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR4_CONTROL(PF0_SRIOV_BAR4_CONTROL)
   ,.PF1_SRIOV_BAR4_CONTROL(PF1_SRIOV_BAR4_CONTROL)
   ,.PF2_SRIOV_BAR4_CONTROL(PF2_SRIOV_BAR4_CONTROL)
   ,.PF3_SRIOV_BAR4_CONTROL(PF3_SRIOV_BAR4_CONTROL)
   ,.PF0_SRIOV_BAR4_APERTURE_SIZE(PF0_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR4_APERTURE_SIZE(PF1_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR4_APERTURE_SIZE(PF2_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR4_APERTURE_SIZE(PF3_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR5_CONTROL(PF0_SRIOV_BAR5_CONTROL)
   ,.PF1_SRIOV_BAR5_CONTROL(PF1_SRIOV_BAR5_CONTROL)
   ,.PF2_SRIOV_BAR5_CONTROL(PF2_SRIOV_BAR5_CONTROL)
   ,.PF3_SRIOV_BAR5_CONTROL(PF3_SRIOV_BAR5_CONTROL)
   ,.PF0_SRIOV_BAR5_APERTURE_SIZE(PF0_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR5_APERTURE_SIZE(PF1_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR5_APERTURE_SIZE(PF2_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR5_APERTURE_SIZE(PF3_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF0_TPHR_CAP_NEXTPTR(PF0_TPHR_CAP_NEXTPTR)
   ,.PF1_TPHR_CAP_NEXTPTR(PF1_TPHR_CAP_NEXTPTR)
   ,.PF2_TPHR_CAP_NEXTPTR(PF2_TPHR_CAP_NEXTPTR)
   ,.PF3_TPHR_CAP_NEXTPTR(PF3_TPHR_CAP_NEXTPTR)
   ,.VFG0_TPHR_CAP_NEXTPTR(VFG0_TPHR_CAP_NEXTPTR)
   ,.VFG1_TPHR_CAP_NEXTPTR(VFG1_TPHR_CAP_NEXTPTR)
   ,.VFG2_TPHR_CAP_NEXTPTR(VFG2_TPHR_CAP_NEXTPTR)
   ,.VFG3_TPHR_CAP_NEXTPTR(VFG3_TPHR_CAP_NEXTPTR)
   ,.PF0_TPHR_CAP_VER(PF0_TPHR_CAP_VER)
   ,.PF0_TPHR_CAP_INT_VEC_MODE(PF0_TPHR_CAP_INT_VEC_MODE)
   ,.PF0_TPHR_CAP_DEV_SPECIFIC_MODE(PF0_TPHR_CAP_DEV_SPECIFIC_MODE)
   ,.PF0_TPHR_CAP_ST_TABLE_LOC(PF0_TPHR_CAP_ST_TABLE_LOC)
   ,.PF0_TPHR_CAP_ST_TABLE_SIZE(PF0_TPHR_CAP_ST_TABLE_SIZE)
   ,.PF0_TPHR_CAP_ST_MODE_SEL(PF0_TPHR_CAP_ST_MODE_SEL)
   ,.PF1_TPHR_CAP_ST_MODE_SEL(PF1_TPHR_CAP_ST_MODE_SEL)
   ,.PF2_TPHR_CAP_ST_MODE_SEL(PF2_TPHR_CAP_ST_MODE_SEL)
   ,.PF3_TPHR_CAP_ST_MODE_SEL(PF3_TPHR_CAP_ST_MODE_SEL)
   ,.VFG0_TPHR_CAP_ST_MODE_SEL(VFG0_TPHR_CAP_ST_MODE_SEL)
   ,.VFG1_TPHR_CAP_ST_MODE_SEL(VFG1_TPHR_CAP_ST_MODE_SEL)
   ,.VFG2_TPHR_CAP_ST_MODE_SEL(VFG2_TPHR_CAP_ST_MODE_SEL)
   ,.VFG3_TPHR_CAP_ST_MODE_SEL(VFG3_TPHR_CAP_ST_MODE_SEL)
   ,.PF0_TPHR_CAP_ENABLE(PF0_TPHR_CAP_ENABLE)
   ,.TPH_TO_RAM_PIPELINE(TPH_TO_RAM_PIPELINE)
   ,.TPH_FROM_RAM_PIPELINE(TPH_FROM_RAM_PIPELINE)
   ,.MCAP_ENABLE(MCAP_ENABLE)
   ,.MCAP_CONFIGURE_OVERRIDE(MCAP_CONFIGURE_OVERRIDE)
   ,.MCAP_CAP_NEXTPTR(MCAP_CAP_NEXTPTR)
   ,.MCAP_VSEC_ID(MCAP_VSEC_ID)
   ,.MCAP_VSEC_REV(MCAP_VSEC_REV)
   ,.MCAP_VSEC_LEN(MCAP_VSEC_LEN)
   ,.MCAP_FPGA_BITSTREAM_VERSION(MCAP_FPGA_BITSTREAM_VERSION)
   ,.MCAP_INTERRUPT_ON_MCAP_EOS(MCAP_INTERRUPT_ON_MCAP_EOS)
   ,.MCAP_INTERRUPT_ON_MCAP_ERROR(MCAP_INTERRUPT_ON_MCAP_ERROR)
   ,.MCAP_INPUT_GATE_DESIGN_SWITCH(MCAP_INPUT_GATE_DESIGN_SWITCH)
   ,.MCAP_EOS_DESIGN_SWITCH(MCAP_EOS_DESIGN_SWITCH)
   ,.MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH(MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH)
   ,.MCAP_GATE_IO_ENABLE_DESIGN_SWITCH(MCAP_GATE_IO_ENABLE_DESIGN_SWITCH)
   ,.SIM_JTAG_IDCODE(SIM_JTAG_IDCODE)
   ,.DEBUG_AXIST_DISABLE_FEATURE_BIT(DEBUG_AXIST_DISABLE_FEATURE_BIT)
   ,.DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS(DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS)
   ,.DEBUG_TL_DISABLE_FC_TIMEOUT(DEBUG_TL_DISABLE_FC_TIMEOUT)
   ,.DEBUG_PL_DISABLE_SCRAMBLING(DEBUG_PL_DISABLE_SCRAMBLING)
   ,.DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL (DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL )
   ,.DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW (DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW )
   ,.DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR(DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR)
   ,.DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR(DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR)
   ,.DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR(DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR)
   ,.DEBUG_PL_SIM_RESET_LFSR(DEBUG_PL_SIM_RESET_LFSR)
   ,.DEBUG_PL_SPARE(DEBUG_PL_SPARE)
   ,.DEBUG_LL_SPARE(DEBUG_LL_SPARE)
   ,.DEBUG_TL_SPARE(DEBUG_TL_SPARE)
   ,.DEBUG_AXI4ST_SPARE(DEBUG_AXI4ST_SPARE)
   ,.DEBUG_CFG_SPARE(DEBUG_CFG_SPARE)
   ,.DEBUG_CAR_SPARE(DEBUG_CAR_SPARE)
   ,.TEST_MODE_PIN_CHAR(TEST_MODE_PIN_CHAR)
   ,.SPARE_BIT0(SPARE_BIT0)
   ,.SPARE_BIT1(SPARE_BIT1)
   ,.SPARE_BIT2(SPARE_BIT2)
   ,.SPARE_BIT3(SPARE_BIT3)
   ,.SPARE_BIT4(SPARE_BIT4)
   ,.SPARE_BIT5(SPARE_BIT5)
   ,.SPARE_BIT6(SPARE_BIT6)
   ,.SPARE_BIT7(SPARE_BIT7)
   ,.SPARE_BIT8(SPARE_BIT8)
   ,.SPARE_BYTE0(SPARE_BYTE0)
   ,.SPARE_BYTE1(SPARE_BYTE1)
   ,.SPARE_BYTE2(SPARE_BYTE2)
   ,.SPARE_BYTE3(SPARE_BYTE3)
   ,.SPARE_WORD0(SPARE_WORD0)
   ,.SPARE_WORD1(SPARE_WORD1)
   ,.SPARE_WORD2(SPARE_WORD2)
   ,.SPARE_WORD3(SPARE_WORD3)

  ) pcie_4_0_pipe_smsw_inst ( 

    .pipe_rx00_char_is_k(pipe_rx00_char_is_k[1:0])
   ,.pipe_rx01_char_is_k(pipe_rx01_char_is_k[1:0])
   ,.pipe_rx02_char_is_k(pipe_rx02_char_is_k[1:0])
   ,.pipe_rx03_char_is_k(pipe_rx03_char_is_k[1:0])
   ,.pipe_rx04_char_is_k(pipe_rx04_char_is_k[1:0])
   ,.pipe_rx05_char_is_k(pipe_rx05_char_is_k[1:0])
   ,.pipe_rx06_char_is_k(pipe_rx06_char_is_k[1:0])
   ,.pipe_rx07_char_is_k(pipe_rx07_char_is_k[1:0])
   ,.pipe_rx08_char_is_k(pipe_rx08_char_is_k[1:0])
   ,.pipe_rx09_char_is_k(pipe_rx09_char_is_k[1:0])
   ,.pipe_rx10_char_is_k(pipe_rx10_char_is_k[1:0])
   ,.pipe_rx11_char_is_k(pipe_rx11_char_is_k[1:0])
   ,.pipe_rx12_char_is_k(pipe_rx12_char_is_k[1:0])
   ,.pipe_rx13_char_is_k(pipe_rx13_char_is_k[1:0])
   ,.pipe_rx14_char_is_k(pipe_rx14_char_is_k[1:0])
   ,.pipe_rx15_char_is_k(pipe_rx15_char_is_k[1:0])
   ,.pipe_rx00_valid(pipe_rx00_valid)
   ,.pipe_rx01_valid(pipe_rx01_valid)
   ,.pipe_rx02_valid(pipe_rx02_valid)
   ,.pipe_rx03_valid(pipe_rx03_valid)
   ,.pipe_rx04_valid(pipe_rx04_valid)
   ,.pipe_rx05_valid(pipe_rx05_valid)
   ,.pipe_rx06_valid(pipe_rx06_valid)
   ,.pipe_rx07_valid(pipe_rx07_valid)
   ,.pipe_rx08_valid(pipe_rx08_valid)
   ,.pipe_rx09_valid(pipe_rx09_valid)
   ,.pipe_rx10_valid(pipe_rx10_valid)
   ,.pipe_rx11_valid(pipe_rx11_valid)
   ,.pipe_rx12_valid(pipe_rx12_valid)
   ,.pipe_rx13_valid(pipe_rx13_valid)
   ,.pipe_rx14_valid(pipe_rx14_valid)
   ,.pipe_rx15_valid(pipe_rx15_valid)
   ,.pipe_rx00_data(pipe_rx00_data[31:0])
   ,.pipe_rx01_data(pipe_rx01_data[31:0])
   ,.pipe_rx02_data(pipe_rx02_data[31:0])
   ,.pipe_rx03_data(pipe_rx03_data[31:0])
   ,.pipe_rx04_data(pipe_rx04_data[31:0])
   ,.pipe_rx05_data(pipe_rx05_data[31:0])
   ,.pipe_rx06_data(pipe_rx06_data[31:0])
   ,.pipe_rx07_data(pipe_rx07_data[31:0])
   ,.pipe_rx08_data( pipe_tx_rate==2'b11 ? pipe_rx00_data[63:32] : pipe_rx08_data[31:0] )
   ,.pipe_rx09_data( pipe_tx_rate==2'b11 ? pipe_rx01_data[63:32] : pipe_rx09_data[31:0] )
   ,.pipe_rx10_data( pipe_tx_rate==2'b11 ? pipe_rx02_data[63:32] : pipe_rx10_data[31:0] )
   ,.pipe_rx11_data( pipe_tx_rate==2'b11 ? pipe_rx03_data[63:32] : pipe_rx11_data[31:0] )
   ,.pipe_rx12_data( pipe_tx_rate==2'b11 ? pipe_rx04_data[63:32] : pipe_rx12_data[31:0] )
   ,.pipe_rx13_data( pipe_tx_rate==2'b11 ? pipe_rx05_data[63:32] : pipe_rx13_data[31:0] )
   ,.pipe_rx14_data( pipe_tx_rate==2'b11 ? pipe_rx06_data[63:32] : pipe_rx14_data[31:0] )
   ,.pipe_rx15_data( pipe_tx_rate==2'b11 ? pipe_rx07_data[63:32] : pipe_rx15_data[31:0] )
   ,.pipe_rx00_polarity(pipe_rx00_polarity)
   ,.pipe_rx01_polarity(pipe_rx01_polarity)
   ,.pipe_rx02_polarity(pipe_rx02_polarity)
   ,.pipe_rx03_polarity(pipe_rx03_polarity)
   ,.pipe_rx04_polarity(pipe_rx04_polarity)
   ,.pipe_rx05_polarity(pipe_rx05_polarity)
   ,.pipe_rx06_polarity(pipe_rx06_polarity)
   ,.pipe_rx07_polarity(pipe_rx07_polarity)
   ,.pipe_rx08_polarity(pipe_rx08_polarity)
   ,.pipe_rx09_polarity(pipe_rx09_polarity)
   ,.pipe_rx10_polarity(pipe_rx10_polarity)
   ,.pipe_rx11_polarity(pipe_rx11_polarity)
   ,.pipe_rx12_polarity(pipe_rx12_polarity)
   ,.pipe_rx13_polarity(pipe_rx13_polarity)
   ,.pipe_rx14_polarity(pipe_rx14_polarity)
   ,.pipe_rx15_polarity(pipe_rx15_polarity)
   ,.pipe_rx00_status(pipe_rx00_status[2:0])
   ,.pipe_rx01_status(pipe_rx01_status[2:0])
   ,.pipe_rx02_status(pipe_rx02_status[2:0])
   ,.pipe_rx03_status(pipe_rx03_status[2:0])
   ,.pipe_rx04_status(pipe_rx04_status[2:0])
   ,.pipe_rx05_status(pipe_rx05_status[2:0])
   ,.pipe_rx06_status(pipe_rx06_status[2:0])
   ,.pipe_rx07_status(pipe_rx07_status[2:0])
   ,.pipe_rx08_status(pipe_rx08_status[2:0])
   ,.pipe_rx09_status(pipe_rx09_status[2:0])
   ,.pipe_rx10_status(pipe_rx10_status[2:0])
   ,.pipe_rx11_status(pipe_rx11_status[2:0])
   ,.pipe_rx12_status(pipe_rx12_status[2:0])
   ,.pipe_rx13_status(pipe_rx13_status[2:0])
   ,.pipe_rx14_status(pipe_rx14_status[2:0])
   ,.pipe_rx15_status(pipe_rx15_status[2:0])
   ,.pipe_rx00_phy_status(pipe_rx00_phy_status)
   ,.pipe_rx01_phy_status(pipe_rx01_phy_status)
   ,.pipe_rx02_phy_status(pipe_rx02_phy_status)
   ,.pipe_rx03_phy_status(pipe_rx03_phy_status)
   ,.pipe_rx04_phy_status(pipe_rx04_phy_status)
   ,.pipe_rx05_phy_status(pipe_rx05_phy_status)
   ,.pipe_rx06_phy_status(pipe_rx06_phy_status)
   ,.pipe_rx07_phy_status(pipe_rx07_phy_status)
   ,.pipe_rx08_phy_status(pipe_rx08_phy_status)
   ,.pipe_rx09_phy_status(pipe_rx09_phy_status)
   ,.pipe_rx10_phy_status(pipe_rx10_phy_status)
   ,.pipe_rx11_phy_status(pipe_rx11_phy_status)
   ,.pipe_rx12_phy_status(pipe_rx12_phy_status)
   ,.pipe_rx13_phy_status(pipe_rx13_phy_status)
   ,.pipe_rx14_phy_status(pipe_rx14_phy_status)
   ,.pipe_rx15_phy_status(pipe_rx15_phy_status)
   ,.pipe_rx00_elec_idle(pipe_rx00_elec_idle)
   ,.pipe_rx01_elec_idle(pipe_rx01_elec_idle)
   ,.pipe_rx02_elec_idle(pipe_rx02_elec_idle)
   ,.pipe_rx03_elec_idle(pipe_rx03_elec_idle)
   ,.pipe_rx04_elec_idle(pipe_rx04_elec_idle)
   ,.pipe_rx05_elec_idle(pipe_rx05_elec_idle)
   ,.pipe_rx06_elec_idle(pipe_rx06_elec_idle)
   ,.pipe_rx07_elec_idle(pipe_rx07_elec_idle)
   ,.pipe_rx08_elec_idle(pipe_rx08_elec_idle)
   ,.pipe_rx09_elec_idle(pipe_rx09_elec_idle)
   ,.pipe_rx10_elec_idle(pipe_rx10_elec_idle)
   ,.pipe_rx11_elec_idle(pipe_rx11_elec_idle)
   ,.pipe_rx12_elec_idle(pipe_rx12_elec_idle)
   ,.pipe_rx13_elec_idle(pipe_rx13_elec_idle)
   ,.pipe_rx14_elec_idle(pipe_rx14_elec_idle)
   ,.pipe_rx15_elec_idle(pipe_rx15_elec_idle)
   ,.pipe_rx00_data_valid(pipe_rx00_data_valid)
   ,.pipe_rx01_data_valid(pipe_rx01_data_valid)
   ,.pipe_rx02_data_valid(pipe_rx02_data_valid)
   ,.pipe_rx03_data_valid(pipe_rx03_data_valid)
   ,.pipe_rx04_data_valid(pipe_rx04_data_valid)
   ,.pipe_rx05_data_valid(pipe_rx05_data_valid)
   ,.pipe_rx06_data_valid(pipe_rx06_data_valid)
   ,.pipe_rx07_data_valid(pipe_rx07_data_valid)
   ,.pipe_rx08_data_valid(pipe_rx08_data_valid)
   ,.pipe_rx09_data_valid(pipe_rx09_data_valid)
   ,.pipe_rx10_data_valid(pipe_rx10_data_valid)
   ,.pipe_rx11_data_valid(pipe_rx11_data_valid)
   ,.pipe_rx12_data_valid(pipe_rx12_data_valid)
   ,.pipe_rx13_data_valid(pipe_rx13_data_valid)
   ,.pipe_rx14_data_valid(pipe_rx14_data_valid)
   ,.pipe_rx15_data_valid(pipe_rx15_data_valid)
   ,.pipe_rx00_start_block(pipe_rx00_start_block[1:0])
   ,.pipe_rx01_start_block(pipe_rx01_start_block[1:0])
   ,.pipe_rx02_start_block(pipe_rx02_start_block[1:0])
   ,.pipe_rx03_start_block(pipe_rx03_start_block[1:0])
   ,.pipe_rx04_start_block(pipe_rx04_start_block[1:0])
   ,.pipe_rx05_start_block(pipe_rx05_start_block[1:0])
   ,.pipe_rx06_start_block(pipe_rx06_start_block[1:0])
   ,.pipe_rx07_start_block(pipe_rx07_start_block[1:0])
   ,.pipe_rx08_start_block(pipe_rx08_start_block[1:0])
   ,.pipe_rx09_start_block(pipe_rx09_start_block[1:0])
   ,.pipe_rx10_start_block(pipe_rx10_start_block[1:0])
   ,.pipe_rx11_start_block(pipe_rx11_start_block[1:0])
   ,.pipe_rx12_start_block(pipe_rx12_start_block[1:0])
   ,.pipe_rx13_start_block(pipe_rx13_start_block[1:0])
   ,.pipe_rx14_start_block(pipe_rx14_start_block[1:0])
   ,.pipe_rx15_start_block(pipe_rx15_start_block[1:0])
   ,.pipe_rx00_sync_header(pipe_rx00_sync_header[1:0])
   ,.pipe_rx01_sync_header(pipe_rx01_sync_header[1:0])
   ,.pipe_rx02_sync_header(pipe_rx02_sync_header[1:0])
   ,.pipe_rx03_sync_header(pipe_rx03_sync_header[1:0])
   ,.pipe_rx04_sync_header(pipe_rx04_sync_header[1:0])
   ,.pipe_rx05_sync_header(pipe_rx05_sync_header[1:0])
   ,.pipe_rx06_sync_header(pipe_rx06_sync_header[1:0])
   ,.pipe_rx07_sync_header(pipe_rx07_sync_header[1:0])
   ,.pipe_rx08_sync_header(pipe_rx08_sync_header[1:0])
   ,.pipe_rx09_sync_header(pipe_rx09_sync_header[1:0])
   ,.pipe_rx10_sync_header(pipe_rx10_sync_header[1:0])
   ,.pipe_rx11_sync_header(pipe_rx11_sync_header[1:0])
   ,.pipe_rx12_sync_header(pipe_rx12_sync_header[1:0])
   ,.pipe_rx13_sync_header(pipe_rx13_sync_header[1:0])
   ,.pipe_rx14_sync_header(pipe_rx14_sync_header[1:0])
   ,.pipe_rx15_sync_header(pipe_rx15_sync_header[1:0])
   ,.pipe_tx00_compliance(pipe_tx00_compliance)
   ,.pipe_tx01_compliance(pipe_tx01_compliance)
   ,.pipe_tx02_compliance(pipe_tx02_compliance)
   ,.pipe_tx03_compliance(pipe_tx03_compliance)
   ,.pipe_tx04_compliance(pipe_tx04_compliance)
   ,.pipe_tx05_compliance(pipe_tx05_compliance)
   ,.pipe_tx06_compliance(pipe_tx06_compliance)
   ,.pipe_tx07_compliance(pipe_tx07_compliance)
   ,.pipe_tx08_compliance(pipe_tx08_compliance)
   ,.pipe_tx09_compliance(pipe_tx09_compliance)
   ,.pipe_tx10_compliance(pipe_tx10_compliance)
   ,.pipe_tx11_compliance(pipe_tx11_compliance)
   ,.pipe_tx12_compliance(pipe_tx12_compliance)
   ,.pipe_tx13_compliance(pipe_tx13_compliance)
   ,.pipe_tx14_compliance(pipe_tx14_compliance)
   ,.pipe_tx15_compliance(pipe_tx15_compliance)
   ,.pipe_tx00_char_is_k(pipe_tx00_char_is_k[1:0])
   ,.pipe_tx01_char_is_k(pipe_tx01_char_is_k[1:0])
   ,.pipe_tx02_char_is_k(pipe_tx02_char_is_k[1:0])
   ,.pipe_tx03_char_is_k(pipe_tx03_char_is_k[1:0])
   ,.pipe_tx04_char_is_k(pipe_tx04_char_is_k[1:0])
   ,.pipe_tx05_char_is_k(pipe_tx05_char_is_k[1:0])
   ,.pipe_tx06_char_is_k(pipe_tx06_char_is_k[1:0])
   ,.pipe_tx07_char_is_k(pipe_tx07_char_is_k[1:0])
   ,.pipe_tx08_char_is_k(pipe_tx08_char_is_k[1:0])
   ,.pipe_tx09_char_is_k(pipe_tx09_char_is_k[1:0])
   ,.pipe_tx10_char_is_k(pipe_tx10_char_is_k[1:0])
   ,.pipe_tx11_char_is_k(pipe_tx11_char_is_k[1:0])
   ,.pipe_tx12_char_is_k(pipe_tx12_char_is_k[1:0])
   ,.pipe_tx13_char_is_k(pipe_tx13_char_is_k[1:0])
   ,.pipe_tx14_char_is_k(pipe_tx14_char_is_k[1:0])
   ,.pipe_tx15_char_is_k(pipe_tx15_char_is_k[1:0])
   ,.pipe_tx00_data(pipe_tx00_data[31:0])
   ,.pipe_tx01_data(pipe_tx01_data[31:0])
   ,.pipe_tx02_data(pipe_tx02_data[31:0])
   ,.pipe_tx03_data(pipe_tx03_data[31:0])
   ,.pipe_tx04_data(pipe_tx04_data[31:0])
   ,.pipe_tx05_data(pipe_tx05_data[31:0])
   ,.pipe_tx06_data(pipe_tx06_data[31:0])
   ,.pipe_tx07_data(pipe_tx07_data[31:0])
   ,.pipe_tx08_data(pipe_tx08_data[31:0])
   ,.pipe_tx09_data(pipe_tx09_data[31:0])
   ,.pipe_tx10_data(pipe_tx10_data[31:0])
   ,.pipe_tx11_data(pipe_tx11_data[31:0])
   ,.pipe_tx12_data(pipe_tx12_data[31:0])
   ,.pipe_tx13_data(pipe_tx13_data[31:0])
   ,.pipe_tx14_data(pipe_tx14_data[31:0])
   ,.pipe_tx15_data(pipe_tx15_data[31:0])
   ,.pipe_tx00_elec_idle(pipe_tx00_elec_idle)
   ,.pipe_tx01_elec_idle(pipe_tx01_elec_idle)
   ,.pipe_tx02_elec_idle(pipe_tx02_elec_idle)
   ,.pipe_tx03_elec_idle(pipe_tx03_elec_idle)
   ,.pipe_tx04_elec_idle(pipe_tx04_elec_idle)
   ,.pipe_tx05_elec_idle(pipe_tx05_elec_idle)
   ,.pipe_tx06_elec_idle(pipe_tx06_elec_idle)
   ,.pipe_tx07_elec_idle(pipe_tx07_elec_idle)
   ,.pipe_tx08_elec_idle(pipe_tx08_elec_idle)
   ,.pipe_tx09_elec_idle(pipe_tx09_elec_idle)
   ,.pipe_tx10_elec_idle(pipe_tx10_elec_idle)
   ,.pipe_tx11_elec_idle(pipe_tx11_elec_idle)
   ,.pipe_tx12_elec_idle(pipe_tx12_elec_idle)
   ,.pipe_tx13_elec_idle(pipe_tx13_elec_idle)
   ,.pipe_tx14_elec_idle(pipe_tx14_elec_idle)
   ,.pipe_tx15_elec_idle(pipe_tx15_elec_idle)
   ,.pipe_tx00_powerdown(pipe_tx00_powerdown[1:0])
   ,.pipe_tx01_powerdown(pipe_tx01_powerdown[1:0])
   ,.pipe_tx02_powerdown(pipe_tx02_powerdown[1:0])
   ,.pipe_tx03_powerdown(pipe_tx03_powerdown[1:0])
   ,.pipe_tx04_powerdown(pipe_tx04_powerdown[1:0])
   ,.pipe_tx05_powerdown(pipe_tx05_powerdown[1:0])
   ,.pipe_tx06_powerdown(pipe_tx06_powerdown[1:0])
   ,.pipe_tx07_powerdown(pipe_tx07_powerdown[1:0])
   ,.pipe_tx08_powerdown(pipe_tx08_powerdown[1:0])
   ,.pipe_tx09_powerdown(pipe_tx09_powerdown[1:0])
   ,.pipe_tx10_powerdown(pipe_tx10_powerdown[1:0])
   ,.pipe_tx11_powerdown(pipe_tx11_powerdown[1:0])
   ,.pipe_tx12_powerdown(pipe_tx12_powerdown[1:0])
   ,.pipe_tx13_powerdown(pipe_tx13_powerdown[1:0])
   ,.pipe_tx14_powerdown(pipe_tx14_powerdown[1:0])
   ,.pipe_tx15_powerdown(pipe_tx15_powerdown[1:0])
   ,.pipe_tx00_data_valid(pipe_tx00_data_valid)
   ,.pipe_tx01_data_valid(pipe_tx01_data_valid)
   ,.pipe_tx02_data_valid(pipe_tx02_data_valid)
   ,.pipe_tx03_data_valid(pipe_tx03_data_valid)
   ,.pipe_tx04_data_valid(pipe_tx04_data_valid)
   ,.pipe_tx05_data_valid(pipe_tx05_data_valid)
   ,.pipe_tx06_data_valid(pipe_tx06_data_valid)
   ,.pipe_tx07_data_valid(pipe_tx07_data_valid)
   ,.pipe_tx08_data_valid(pipe_tx08_data_valid)
   ,.pipe_tx09_data_valid(pipe_tx09_data_valid)
   ,.pipe_tx10_data_valid(pipe_tx10_data_valid)
   ,.pipe_tx11_data_valid(pipe_tx11_data_valid)
   ,.pipe_tx12_data_valid(pipe_tx12_data_valid)
   ,.pipe_tx13_data_valid(pipe_tx13_data_valid)
   ,.pipe_tx14_data_valid(pipe_tx14_data_valid)
   ,.pipe_tx15_data_valid(pipe_tx15_data_valid)
   ,.pipe_tx00_start_block(pipe_tx00_start_block)
   ,.pipe_tx01_start_block(pipe_tx01_start_block)
   ,.pipe_tx02_start_block(pipe_tx02_start_block)
   ,.pipe_tx03_start_block(pipe_tx03_start_block)
   ,.pipe_tx04_start_block(pipe_tx04_start_block)
   ,.pipe_tx05_start_block(pipe_tx05_start_block)
   ,.pipe_tx06_start_block(pipe_tx06_start_block)
   ,.pipe_tx07_start_block(pipe_tx07_start_block)
   ,.pipe_tx08_start_block(pipe_tx08_start_block)
   ,.pipe_tx09_start_block(pipe_tx09_start_block)
   ,.pipe_tx10_start_block(pipe_tx10_start_block)
   ,.pipe_tx11_start_block(pipe_tx11_start_block)
   ,.pipe_tx12_start_block(pipe_tx12_start_block)
   ,.pipe_tx13_start_block(pipe_tx13_start_block)
   ,.pipe_tx14_start_block(pipe_tx14_start_block)
   ,.pipe_tx15_start_block(pipe_tx15_start_block)
   ,.pipe_tx00_sync_header(pipe_tx00_sync_header[1:0])
   ,.pipe_tx01_sync_header(pipe_tx01_sync_header[1:0])
   ,.pipe_tx02_sync_header(pipe_tx02_sync_header[1:0])
   ,.pipe_tx03_sync_header(pipe_tx03_sync_header[1:0])
   ,.pipe_tx04_sync_header(pipe_tx04_sync_header[1:0])
   ,.pipe_tx05_sync_header(pipe_tx05_sync_header[1:0])
   ,.pipe_tx06_sync_header(pipe_tx06_sync_header[1:0])
   ,.pipe_tx07_sync_header(pipe_tx07_sync_header[1:0])
   ,.pipe_tx08_sync_header(pipe_tx08_sync_header[1:0])
   ,.pipe_tx09_sync_header(pipe_tx09_sync_header[1:0])
   ,.pipe_tx10_sync_header(pipe_tx10_sync_header[1:0])
   ,.pipe_tx11_sync_header(pipe_tx11_sync_header[1:0])
   ,.pipe_tx12_sync_header(pipe_tx12_sync_header[1:0])
   ,.pipe_tx13_sync_header(pipe_tx13_sync_header[1:0])
   ,.pipe_tx14_sync_header(pipe_tx14_sync_header[1:0])
   ,.pipe_tx15_sync_header(pipe_tx15_sync_header[1:0])
   ,.pipe_rx00_eq_control(pipe_rx00_eq_control[1:0])
   ,.pipe_rx01_eq_control(pipe_rx01_eq_control[1:0])
   ,.pipe_rx02_eq_control(pipe_rx02_eq_control[1:0])
   ,.pipe_rx03_eq_control(pipe_rx03_eq_control[1:0])
   ,.pipe_rx04_eq_control(pipe_rx04_eq_control[1:0])
   ,.pipe_rx05_eq_control(pipe_rx05_eq_control[1:0])
   ,.pipe_rx06_eq_control(pipe_rx06_eq_control[1:0])
   ,.pipe_rx07_eq_control(pipe_rx07_eq_control[1:0])
   ,.pipe_rx08_eq_control(pipe_rx08_eq_control[1:0])
   ,.pipe_rx09_eq_control(pipe_rx09_eq_control[1:0])
   ,.pipe_rx10_eq_control(pipe_rx10_eq_control[1:0])
   ,.pipe_rx11_eq_control(pipe_rx11_eq_control[1:0])
   ,.pipe_rx12_eq_control(pipe_rx12_eq_control[1:0])
   ,.pipe_rx13_eq_control(pipe_rx13_eq_control[1:0])
   ,.pipe_rx14_eq_control(pipe_rx14_eq_control[1:0])
   ,.pipe_rx15_eq_control(pipe_rx15_eq_control[1:0])
   ,.pipe_rx00_eq_lp_lf_fs_sel(pipe_rx00_eq_lp_lf_fs_sel)
   ,.pipe_rx01_eq_lp_lf_fs_sel(pipe_rx01_eq_lp_lf_fs_sel)
   ,.pipe_rx02_eq_lp_lf_fs_sel(pipe_rx02_eq_lp_lf_fs_sel)
   ,.pipe_rx03_eq_lp_lf_fs_sel(pipe_rx03_eq_lp_lf_fs_sel)
   ,.pipe_rx04_eq_lp_lf_fs_sel(pipe_rx04_eq_lp_lf_fs_sel)
   ,.pipe_rx05_eq_lp_lf_fs_sel(pipe_rx05_eq_lp_lf_fs_sel)
   ,.pipe_rx06_eq_lp_lf_fs_sel(pipe_rx06_eq_lp_lf_fs_sel)
   ,.pipe_rx07_eq_lp_lf_fs_sel(pipe_rx07_eq_lp_lf_fs_sel)
   ,.pipe_rx08_eq_lp_lf_fs_sel(pipe_rx08_eq_lp_lf_fs_sel)
   ,.pipe_rx09_eq_lp_lf_fs_sel(pipe_rx09_eq_lp_lf_fs_sel)
   ,.pipe_rx10_eq_lp_lf_fs_sel(pipe_rx10_eq_lp_lf_fs_sel)
   ,.pipe_rx11_eq_lp_lf_fs_sel(pipe_rx11_eq_lp_lf_fs_sel)
   ,.pipe_rx12_eq_lp_lf_fs_sel(pipe_rx12_eq_lp_lf_fs_sel)
   ,.pipe_rx13_eq_lp_lf_fs_sel(pipe_rx13_eq_lp_lf_fs_sel)
   ,.pipe_rx14_eq_lp_lf_fs_sel(pipe_rx14_eq_lp_lf_fs_sel)
   ,.pipe_rx15_eq_lp_lf_fs_sel(pipe_rx15_eq_lp_lf_fs_sel)
   ,.pipe_rx00_eq_lp_new_tx_coeff_or_preset(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx01_eq_lp_new_tx_coeff_or_preset(pipe_rx01_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx02_eq_lp_new_tx_coeff_or_preset(pipe_rx02_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx03_eq_lp_new_tx_coeff_or_preset(pipe_rx03_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx04_eq_lp_new_tx_coeff_or_preset(pipe_rx04_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx05_eq_lp_new_tx_coeff_or_preset(pipe_rx05_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx06_eq_lp_new_tx_coeff_or_preset(pipe_rx06_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx07_eq_lp_new_tx_coeff_or_preset(pipe_rx07_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx08_eq_lp_new_tx_coeff_or_preset(pipe_rx08_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx09_eq_lp_new_tx_coeff_or_preset(pipe_rx09_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx10_eq_lp_new_tx_coeff_or_preset(pipe_rx10_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx11_eq_lp_new_tx_coeff_or_preset(pipe_rx11_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx12_eq_lp_new_tx_coeff_or_preset(pipe_rx12_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx13_eq_lp_new_tx_coeff_or_preset(pipe_rx13_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx14_eq_lp_new_tx_coeff_or_preset(pipe_rx14_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx15_eq_lp_new_tx_coeff_or_preset(pipe_rx15_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx00_eq_lp_adapt_done(pipe_rx00_eq_lp_adapt_done)
   ,.pipe_rx01_eq_lp_adapt_done(pipe_rx01_eq_lp_adapt_done)
   ,.pipe_rx02_eq_lp_adapt_done(pipe_rx02_eq_lp_adapt_done)
   ,.pipe_rx03_eq_lp_adapt_done(pipe_rx03_eq_lp_adapt_done)
   ,.pipe_rx04_eq_lp_adapt_done(pipe_rx04_eq_lp_adapt_done)
   ,.pipe_rx05_eq_lp_adapt_done(pipe_rx05_eq_lp_adapt_done)
   ,.pipe_rx06_eq_lp_adapt_done(pipe_rx06_eq_lp_adapt_done)
   ,.pipe_rx07_eq_lp_adapt_done(pipe_rx07_eq_lp_adapt_done)
   ,.pipe_rx08_eq_lp_adapt_done(pipe_rx08_eq_lp_adapt_done)
   ,.pipe_rx09_eq_lp_adapt_done(pipe_rx09_eq_lp_adapt_done)
   ,.pipe_rx10_eq_lp_adapt_done(pipe_rx10_eq_lp_adapt_done)
   ,.pipe_rx11_eq_lp_adapt_done(pipe_rx11_eq_lp_adapt_done)
   ,.pipe_rx12_eq_lp_adapt_done(pipe_rx12_eq_lp_adapt_done)
   ,.pipe_rx13_eq_lp_adapt_done(pipe_rx13_eq_lp_adapt_done)
   ,.pipe_rx14_eq_lp_adapt_done(pipe_rx14_eq_lp_adapt_done)
   ,.pipe_rx15_eq_lp_adapt_done(pipe_rx15_eq_lp_adapt_done)
   ,.pipe_rx00_eq_done(pipe_rx00_eq_done)
   ,.pipe_rx01_eq_done(pipe_rx01_eq_done)
   ,.pipe_rx02_eq_done(pipe_rx02_eq_done)
   ,.pipe_rx03_eq_done(pipe_rx03_eq_done)
   ,.pipe_rx04_eq_done(pipe_rx04_eq_done)
   ,.pipe_rx05_eq_done(pipe_rx05_eq_done)
   ,.pipe_rx06_eq_done(pipe_rx06_eq_done)
   ,.pipe_rx07_eq_done(pipe_rx07_eq_done)
   ,.pipe_rx08_eq_done(pipe_rx08_eq_done)
   ,.pipe_rx09_eq_done(pipe_rx09_eq_done)
   ,.pipe_rx10_eq_done(pipe_rx10_eq_done)
   ,.pipe_rx11_eq_done(pipe_rx11_eq_done)
   ,.pipe_rx12_eq_done(pipe_rx12_eq_done)
   ,.pipe_rx13_eq_done(pipe_rx13_eq_done)
   ,.pipe_rx14_eq_done(pipe_rx14_eq_done)
   ,.pipe_rx15_eq_done(pipe_rx15_eq_done)
   ,.pipe_tx00_eq_control(pipe_tx00_eq_control[1:0])
   ,.pipe_tx01_eq_control(pipe_tx01_eq_control[1:0])
   ,.pipe_tx02_eq_control(pipe_tx02_eq_control[1:0])
   ,.pipe_tx03_eq_control(pipe_tx03_eq_control[1:0])
   ,.pipe_tx04_eq_control(pipe_tx04_eq_control[1:0])
   ,.pipe_tx05_eq_control(pipe_tx05_eq_control[1:0])
   ,.pipe_tx06_eq_control(pipe_tx06_eq_control[1:0])
   ,.pipe_tx07_eq_control(pipe_tx07_eq_control[1:0])
   ,.pipe_tx08_eq_control(pipe_tx08_eq_control[1:0])
   ,.pipe_tx09_eq_control(pipe_tx09_eq_control[1:0])
   ,.pipe_tx10_eq_control(pipe_tx10_eq_control[1:0])
   ,.pipe_tx11_eq_control(pipe_tx11_eq_control[1:0])
   ,.pipe_tx12_eq_control(pipe_tx12_eq_control[1:0])
   ,.pipe_tx13_eq_control(pipe_tx13_eq_control[1:0])
   ,.pipe_tx14_eq_control(pipe_tx14_eq_control[1:0])
   ,.pipe_tx15_eq_control(pipe_tx15_eq_control[1:0])
   ,.pipe_tx00_eq_deemph(pipe_tx00_eq_deemph[5:0])
   ,.pipe_tx01_eq_deemph(pipe_tx01_eq_deemph[5:0])
   ,.pipe_tx02_eq_deemph(pipe_tx02_eq_deemph[5:0])
   ,.pipe_tx03_eq_deemph(pipe_tx03_eq_deemph[5:0])
   ,.pipe_tx04_eq_deemph(pipe_tx04_eq_deemph[5:0])
   ,.pipe_tx05_eq_deemph(pipe_tx05_eq_deemph[5:0])
   ,.pipe_tx06_eq_deemph(pipe_tx06_eq_deemph[5:0])
   ,.pipe_tx07_eq_deemph(pipe_tx07_eq_deemph[5:0])
   ,.pipe_tx08_eq_deemph(pipe_tx08_eq_deemph[5:0])
   ,.pipe_tx09_eq_deemph(pipe_tx09_eq_deemph[5:0])
   ,.pipe_tx10_eq_deemph(pipe_tx10_eq_deemph[5:0])
   ,.pipe_tx11_eq_deemph(pipe_tx11_eq_deemph[5:0])
   ,.pipe_tx12_eq_deemph(pipe_tx12_eq_deemph[5:0])
   ,.pipe_tx13_eq_deemph(pipe_tx13_eq_deemph[5:0])
   ,.pipe_tx14_eq_deemph(pipe_tx14_eq_deemph[5:0])
   ,.pipe_tx15_eq_deemph(pipe_tx15_eq_deemph[5:0])
   ,.pipe_tx00_eq_coeff(pipe_tx00_eq_coeff[17:0])
   ,.pipe_tx01_eq_coeff(pipe_tx01_eq_coeff[17:0])
   ,.pipe_tx02_eq_coeff(pipe_tx02_eq_coeff[17:0])
   ,.pipe_tx03_eq_coeff(pipe_tx03_eq_coeff[17:0])
   ,.pipe_tx04_eq_coeff(pipe_tx04_eq_coeff[17:0])
   ,.pipe_tx05_eq_coeff(pipe_tx05_eq_coeff[17:0])
   ,.pipe_tx06_eq_coeff(pipe_tx06_eq_coeff[17:0])
   ,.pipe_tx07_eq_coeff(pipe_tx07_eq_coeff[17:0])
   ,.pipe_tx08_eq_coeff(pipe_tx08_eq_coeff[17:0])
   ,.pipe_tx09_eq_coeff(pipe_tx09_eq_coeff[17:0])
   ,.pipe_tx10_eq_coeff(pipe_tx10_eq_coeff[17:0])
   ,.pipe_tx11_eq_coeff(pipe_tx11_eq_coeff[17:0])
   ,.pipe_tx12_eq_coeff(pipe_tx12_eq_coeff[17:0])
   ,.pipe_tx13_eq_coeff(pipe_tx13_eq_coeff[17:0])
   ,.pipe_tx14_eq_coeff(pipe_tx14_eq_coeff[17:0])
   ,.pipe_tx15_eq_coeff(pipe_tx15_eq_coeff[17:0])
   ,.pipe_tx00_eq_done(pipe_tx00_eq_done)
   ,.pipe_tx01_eq_done(pipe_tx01_eq_done)
   ,.pipe_tx02_eq_done(pipe_tx02_eq_done)
   ,.pipe_tx03_eq_done(pipe_tx03_eq_done)
   ,.pipe_tx04_eq_done(pipe_tx04_eq_done)
   ,.pipe_tx05_eq_done(pipe_tx05_eq_done)
   ,.pipe_tx06_eq_done(pipe_tx06_eq_done)
   ,.pipe_tx07_eq_done(pipe_tx07_eq_done)
   ,.pipe_tx08_eq_done(pipe_tx08_eq_done)
   ,.pipe_tx09_eq_done(pipe_tx09_eq_done)
   ,.pipe_tx10_eq_done(pipe_tx10_eq_done)
   ,.pipe_tx11_eq_done(pipe_tx11_eq_done)
   ,.pipe_tx12_eq_done(pipe_tx12_eq_done)
   ,.pipe_tx13_eq_done(pipe_tx13_eq_done)
   ,.pipe_tx14_eq_done(pipe_tx14_eq_done)
   ,.pipe_tx15_eq_done(pipe_tx15_eq_done)
   ,.pipe_rx_eq_lp_tx_preset(pipe_rx_eq_lp_tx_preset[3:0])
   ,.pipe_rx_eq_lp_lf_fs(pipe_rx_eq_lp_lf_fs[5:0])
   ,.pipe_tx_rcvr_det(pipe_tx_rcvr_det)
   ,.pipe_tx_rate(pipe_tx_rate[1:0])
   ,.pipe_tx_deemph(pipe_tx_deemph)
   ,.pipe_tx_margin(pipe_tx_margin[2:0])
   ,.pipe_tx_swing(pipe_tx_swing)
   ,.pipe_tx_reset(pipe_tx_reset)
   ,.pipe_eq_fs(pipe_eq_fs[5:0])
   ,.pipe_eq_lf(pipe_eq_lf[5:0])
   ,.pl_gen2_upstream_prefer_deemph(pl_gen2_upstream_prefer_deemph)
   ,.pl_eq_in_progress(pl_eq_in_progress)
   ,.pl_eq_phase(pl_eq_phase[1:0])
   ,.pl_eq_reset_eieos_count(1'b0)
   ,.pl_redo_eq(pl_redo_eq)
   ,.pl_redo_eq_speed(pl_redo_eq_speed)
   ,.pl_eq_mismatch(pl_eq_mismatch)
   ,.pl_redo_eq_pending(pl_redo_eq_pending)
   ,.m_axis_cq_tdata(m_axis_cq_tdata[AXI4_DATA_WIDTH-1:0])
   ,.s_axis_cc_tdata(s_axis_cc_tdata[AXI4_DATA_WIDTH-1:0])
   ,.s_axis_rq_tdata(s_axis_rq_tdata[AXI4_DATA_WIDTH-1:0])
   ,.m_axis_rc_tdata(m_axis_rc_tdata[AXI4_DATA_WIDTH-1:0])
   ,.m_axis_cq_tuser(m_axis_cq_tuser[AXI4_CQ_TUSER_WIDTH-1:0])
   ,.s_axis_cc_tuser(s_axis_cc_tuser[AXI4_CC_TUSER_WIDTH-1:0])
   ,.m_axis_cq_tlast(m_axis_cq_tlast)
   ,.s_axis_rq_tlast(s_axis_rq_tlast)
   ,.m_axis_rc_tlast(m_axis_rc_tlast)
   ,.s_axis_cc_tlast(s_axis_cc_tlast)
   ,.pcie_cq_np_req(pcie_cq_np_req[1:0])
   ,.pcie_cq_np_req_count(pcie_cq_np_req_count[5:0])
   ,.s_axis_rq_tuser(s_axis_rq_tuser[AXI4_RQ_TUSER_WIDTH-1:0])
   ,.m_axis_rc_tuser(m_axis_rc_tuser[AXI4_RC_TUSER_WIDTH-1:0])
   ,.m_axis_cq_tkeep(m_axis_cq_tkeep[AXI4_TKEEP_WIDTH-1:0])
   ,.s_axis_cc_tkeep(s_axis_cc_tkeep[AXI4_TKEEP_WIDTH-1:0])
   ,.s_axis_rq_tkeep(s_axis_rq_tkeep[AXI4_TKEEP_WIDTH-1:0])
   ,.m_axis_rc_tkeep(m_axis_rc_tkeep[AXI4_TKEEP_WIDTH-1:0])
   ,.m_axis_cq_tvalid(m_axis_cq_tvalid)
   ,.s_axis_cc_tvalid(s_axis_cc_tvalid)
   ,.s_axis_rq_tvalid(s_axis_rq_tvalid)
   ,.m_axis_rc_tvalid(m_axis_rc_tvalid)
   ,.m_axis_cq_tready({AXI4_CQ_TREADY_WIDTH{m_axis_cq_tready}})
   ,.s_axis_cc_tready(s_axis_cc_tready)
   ,.s_axis_rq_tready(s_axis_rq_tready)
   ,.m_axis_rc_tready({AXI4_RC_TREADY_WIDTH{m_axis_rc_tready}})
   ,.pcie_rq_seq_num0(pcie_rq_seq_num0[5:0])
   ,.pcie_rq_seq_num_vld0(pcie_rq_seq_num_vld0)
   ,.pcie_rq_seq_num1(pcie_rq_seq_num1[5:0])
   ,.pcie_rq_seq_num_vld1(pcie_rq_seq_num_vld1)
   ,.pcie_rq_tag0(pcie_rq_tag0[7:0])
   ,.pcie_rq_tag_vld0(pcie_rq_tag_vld0)
   ,.pcie_rq_tag1(pcie_rq_tag1[7:0])
   ,.pcie_rq_tag_vld1(pcie_rq_tag_vld1)
   ,.pcie_tfc_nph_av(pcie_tfc_nph_av[3:0])
   ,.pcie_tfc_npd_av(pcie_tfc_npd_av[3:0])
   ,.pcie_rq_tag_av(pcie_rq_tag_av[3:0])
   ,.axi_user_out( )
   ,.axi_user_in(8'h00)
   ,.cfg_mgmt_addr(cfg_mgmt_addr[9:0])
   ,.cfg_mgmt_function_number(cfg_mgmt_function_number[7:0])
   ,.cfg_mgmt_write(cfg_mgmt_write)
   ,.cfg_mgmt_write_data(cfg_mgmt_write_data[31:0])
   ,.cfg_mgmt_byte_enable(cfg_mgmt_byte_enable[3:0])
   ,.cfg_mgmt_read(cfg_mgmt_read)
   ,.cfg_mgmt_read_data(cfg_mgmt_read_data[31:0])
   ,.cfg_mgmt_read_write_done(cfg_mgmt_read_write_done)
   ,.cfg_mgmt_debug_access(cfg_mgmt_debug_access)
   ,.cfg_phy_link_down(cfg_phy_link_down)
   ,.cfg_phy_link_status(cfg_phy_link_status[1:0])
   ,.cfg_negotiated_width(cfg_negotiated_width[2:0])
   ,.cfg_current_speed(cfg_current_speed[1:0])
   ,.cfg_max_payload(cfg_max_payload[1:0])
   ,.cfg_max_read_req(cfg_max_read_req[2:0])
   ,.cfg_function_status(cfg_function_status[15:0])
   ,.cfg_function_power_state(cfg_function_power_state[11:0])
   ,.cfg_link_power_state(cfg_link_power_state[1:0])
   ,.cfg_err_cor_out(cfg_err_cor_out)
   ,.cfg_err_nonfatal_out(cfg_err_nonfatal_out)
   ,.cfg_err_fatal_out(cfg_err_fatal_out)
   ,.cfg_local_error_valid(cfg_local_error_valid)
   ,.cfg_local_error_out(cfg_local_error_out[4:0])
   ,.cfg_ltr_enable()
   ,.cfg_ltssm_state(cfg_ltssm_state[5:0])
   ,.cfg_rx_pm_state(cfg_rx_pm_state[1:0])
   ,.cfg_tx_pm_state(cfg_tx_pm_state[1:0])
   ,.cfg_rcb_status(cfg_rcb_status[3:0])
   ,.cfg_obff_enable(cfg_obff_enable[1:0])
   ,.cfg_pl_status_change(cfg_pl_status_change)
   ,.cfg_tph_requester_enable(cfg_tph_requester_enable[3:0])
   ,.cfg_tph_st_mode(cfg_tph_st_mode[11:0])
   ,.cfg_msg_received(cfg_msg_received)
   ,.cfg_msg_received_data(cfg_msg_received_data[7:0])
   ,.cfg_msg_received_type(cfg_msg_received_type[4:0])
   ,.cfg_msg_transmit(cfg_msg_transmit_int)
   ,.cfg_msg_transmit_type(cfg_msg_transmit_type[2:0])
   ,.cfg_msg_transmit_data(cfg_msg_transmit_data[31:0])
   ,.cfg_msg_transmit_done(cfg_msg_transmit_done)
   ,.cfg_fc_ph(cfg_fc_ph[7:0])
   ,.cfg_fc_pd(cfg_fc_pd[11:0])
   ,.cfg_fc_nph(cfg_fc_nph[7:0])
   ,.cfg_fc_npd(cfg_fc_npd[11:0])
   ,.cfg_fc_cplh(cfg_fc_cplh[7:0])
   ,.cfg_fc_cpld(cfg_fc_cpld[11:0])
   ,.cfg_fc_sel(cfg_fc_sel[2:0])
   ,.cfg_hot_reset_in(cfg_hot_reset_in)
   ,.cfg_hot_reset_out(cfg_hot_reset_out)
   ,.cfg_config_space_enable(cfg_config_space_enable)
   ,.cfg_dsn(cfg_dsn[63:0])
   ,.cfg_dev_id_pf0(cfg_dev_id_pf0[15:0])
   ,.cfg_dev_id_pf1(cfg_dev_id_pf1[15:0])
   ,.cfg_dev_id_pf2(cfg_dev_id_pf2[15:0])
   ,.cfg_dev_id_pf3(cfg_dev_id_pf3[15:0])
   ,.cfg_vend_id(cfg_vend_id[15:0])
   ,.cfg_rev_id_pf0(cfg_rev_id_pf0[7:0])
   ,.cfg_rev_id_pf1(cfg_rev_id_pf1[7:0])
   ,.cfg_rev_id_pf2(cfg_rev_id_pf2[7:0])
   ,.cfg_rev_id_pf3(cfg_rev_id_pf3[7:0])
   ,.cfg_subsys_id_pf0(cfg_subsys_id_pf0[15:0])
   ,.cfg_subsys_id_pf1(cfg_subsys_id_pf1[15:0])
   ,.cfg_subsys_id_pf2(cfg_subsys_id_pf2[15:0])
   ,.cfg_subsys_id_pf3(cfg_subsys_id_pf3[15:0])
   ,.cfg_subsys_vend_id(cfg_subsys_vend_id[15:0])
   ,.cfg_ds_port_number(cfg_ds_port_number[7:0])
   ,.cfg_ds_bus_number(cfg_ds_bus_number[7:0])
   ,.cfg_ds_device_number(cfg_ds_device_number[4:0])
   ,.cfg_ds_function_number(3'b0)
   ,.cfg_bus_number(cfg_bus_number[7:0])
   ,.cfg_power_state_change_ack(cfg_power_state_change_ack)
   ,.cfg_power_state_change_interrupt(cfg_power_state_change_interrupt)
   ,.cfg_err_cor_in(cfg_err_cor_in)
   ,.cfg_err_uncor_in(cfg_err_uncor_in)
   ,.cfg_flr_done(cfg_flr_done[3:0])
   ,.cfg_vf_flr_in_process(cfg_vf_flr_in_process[251:0])   
   ,.cfg_vf_flr_done(cfg_vf_flr_done)                      
   ,.cfg_vf_flr_func_num(cfg_vf_flr_func_num[7:0])
   ,.cfg_vf_status(cfg_vf_status[503:0])                   
   ,.cfg_vf_power_state(cfg_vf_power_state[755:0])         
   ,.cfg_vf_tph_requester_enable( cfg_vf_tph_requester_enable[251:0])
   ,.cfg_vf_tph_st_mode(cfg_vf_tph_st_mode[755:0])         
   ,.cfg_interrupt_msix_vf_enable(cfg_interrupt_msix_vf_enable[251:0])
   ,.cfg_interrupt_msix_vf_mask(cfg_interrupt_msix_vf_mask[251:0])
   ,.cfg_flr_in_process(cfg_flr_in_process[3:0])
   ,.cfg_req_pm_transition_l23_ready(cfg_req_pm_transition_l23_ready)
   ,.cfg_link_training_enable(cfg_link_training_enable)
   ,.cfg_interrupt_int(cfg_interrupt_int[3:0])
   ,.cfg_interrupt_sent(cfg_interrupt_sent)
   ,.cfg_interrupt_pending(cfg_interrupt_pending[3:0])
   ,.cfg_interrupt_msi_enable(cfg_interrupt_msi_enable[3:0])
   ,.cfg_interrupt_msi_int(cfg_interrupt_msi_int[31:0])
   ,.cfg_interrupt_msi_sent(cfg_interrupt_msi_sent)
   ,.cfg_interrupt_msi_fail(cfg_interrupt_msi_fail)
   ,.cfg_interrupt_msi_mmenable(cfg_interrupt_msi_mmenable[11:0])
   ,.cfg_interrupt_msi_pending_status(cfg_interrupt_msi_pending_status[31:0])
   ,.cfg_interrupt_msi_pending_status_function_num(cfg_interrupt_msi_pending_status_function_num[1:0])
   ,.cfg_interrupt_msi_pending_status_data_enable(cfg_interrupt_msi_pending_status_data_enable)
   ,.cfg_interrupt_msi_mask_update(cfg_interrupt_msi_mask_update)
   ,.cfg_interrupt_msi_select(cfg_interrupt_msi_select[1:0])
   ,.cfg_interrupt_msi_data(cfg_interrupt_msi_data[31:0])
   ,.cfg_interrupt_msix_enable(cfg_interrupt_msix_enable[3:0])
   ,.cfg_interrupt_msix_mask(cfg_interrupt_msix_mask[3:0])
   ,.cfg_interrupt_msix_address(cfg_interrupt_msix_address[63:0])
   ,.cfg_interrupt_msix_data(cfg_interrupt_msix_data[31:0])
   ,.cfg_interrupt_msix_int(cfg_interrupt_msix_int)
   ,.cfg_interrupt_msix_vec_pending(cfg_interrupt_msix_vec_pending[1:0])
   ,.cfg_interrupt_msix_vec_pending_status(cfg_interrupt_msix_vec_pending_status)
   ,.cfg_interrupt_msi_attr(cfg_interrupt_msi_attr[2:0])
   ,.cfg_interrupt_msi_tph_present(cfg_interrupt_msi_tph_present)
   ,.cfg_interrupt_msi_tph_type(cfg_interrupt_msi_tph_type[1:0])
   ,.cfg_interrupt_msi_tph_st_tag(cfg_interrupt_msi_tph_st_tag[7:0])
   ,.cfg_interrupt_msi_function_number(cfg_interrupt_msi_function_number[7:0])
   ,.cfg_ext_read_received(cfg_ext_read_received)
   ,.cfg_ext_write_received(cfg_ext_write_received)
   ,.cfg_ext_register_number(cfg_ext_register_number[9:0])
   ,.cfg_ext_function_number(cfg_ext_function_number[7:0])
   ,.cfg_ext_write_data(cfg_ext_write_data[31:0])
   ,.cfg_ext_write_byte_enable(cfg_ext_write_byte_enable[3:0])
   ,.cfg_ext_read_data(cfg_ext_read_data[31:0])
   ,.cfg_ext_read_data_valid(cfg_ext_read_data_valid)
   ,.cfg_pm_aspm_l1_entry_reject(cfg_pm_aspm_l1_entry_reject)
   ,.cfg_pm_aspm_tx_l0s_entry_disable(cfg_pm_aspm_tx_l0s_entry_disable)
   ,.user_tph_stt_func_num(8'h00)
   ,.user_tph_stt_index(6'b0)
   ,.user_tph_stt_rd_en(1'b0)
   ,.user_tph_stt_rd_data()
   ,.conf_req_type(conf_req_type[1:0])
   ,.conf_req_reg_num(conf_req_reg_num[3:0])
   ,.conf_req_data(conf_req_data[31:0])
   ,.conf_req_valid(conf_req_valid)
   ,.conf_req_ready(conf_req_ready)
   ,.conf_resp_rdata(conf_resp_rdata[31:0])
   ,.conf_resp_valid(conf_resp_valid)
   ,.conf_mcap_design_switch(conf_mcap_design_switch)
   ,.conf_mcap_eos(conf_mcap_eos)
   ,.conf_mcap_in_use_by_pcie(conf_mcap_in_use_by_pcie)
   ,.conf_mcap_request_by_conf(conf_mcap_request_by_conf)

   ,.drp_clk('h0)
   ,.drp_en('h0)
   ,.drp_we('h0)
   ,.drp_addr('h0)
   ,.drp_di('h0)
   ,.drp_rdy()
   ,.drp_do()
   ,.pipe_clk(pipe_clk)
   ,.core_clk(core_clk)
   ,.user_clk(user_clk)
   ,.user_clk2(user_clk2)
   ,.user_clk_en(user_clk_en)
   ,.mcap_clk(mcap_clk)
   ,.mcap_rst_b(mcap_rst_b)
   ,.pcie_perst0_b(pcie_perst0_b)
   ,.pcie_perst1_b(pcie_perst1_b)
   ,.phy_rdy(phy_rdy)

  );

  BUFG_GT bufg_gt_sysclk (.CE (1'd1), .CEMASK (1'd0), .CLR (1'd0), .CLRMASK (1'd0), .DIV (3'd0), .I (sys_clk), .O (sys_clk_bufg));

  always @(posedge user_clk or posedge sys_or_hot_rst) begin
   if (sys_or_hot_rst) begin
      as_cdr_hold_req_user    <= 1'b0;
      as_mac_in_detect_user   <= 1'b1;
   end else begin
      // If LTSSM state is Recovery.Speed, L1.Entry, L1.Idle, Loopback.Entry_slave, or Loopback.Speed
      as_cdr_hold_req_user    <= (cfg_ltssm_state == 6'h0C) | (cfg_ltssm_state == 6'h17) |
                                 (cfg_ltssm_state == 6'h18) | (cfg_ltssm_state == 6'h24) |
                                 (cfg_ltssm_state == 6'h2D);
      // If LTSSM state is Detect.Quiet or Detect.Active
      as_mac_in_detect_user   <= (cfg_ltssm_state == 6'h00) | (cfg_ltssm_state == 6'h01);
   end
  end

  // Sync to PIPE_CLK
  always @(posedge pipe_clk or posedge sys_or_hot_rst) begin
   if (sys_or_hot_rst) begin
      as_cdr_hold_req_ff    <= 1'b0;
      as_cdr_hold_req_ff1   <= 1'b0;
      as_mac_in_detect_ff   <= 1'b1;
      as_mac_in_detect_ff1  <= 1'b1;
   end else begin
      as_cdr_hold_req_ff    <= as_cdr_hold_req_user;
      as_cdr_hold_req_ff1   <= as_cdr_hold_req_ff;
      as_mac_in_detect_ff   <= as_mac_in_detect_user;
      as_mac_in_detect_ff1  <= as_mac_in_detect_ff;
   end
  end

xp4_usp_smsw_phy_top #
  (
    //--------------------------------------------------------------------------
    //  Parameters
    //--------------------------------------------------------------------------
    .FPGA_FAMILY      ( FPGA_FAMILY ),
    .FPGA_XCVR        ( FPGA_XCVR ),
    .PIPELINE_STAGES  ( PIPE_PIPELINE_STAGES ),
    .PHY_SIM_EN       ( ((PL_SIM_FAST_LINK_TRAINING != 2'b0) ? "TRUE" : "FALSE") ),     
    .PHY_LANE         ( PL_LINK_CAP_MAX_LINK_WIDTH ),   
    .PHY_MAX_SPEED    ( (PL_LINK_CAP_MAX_LINK_SPEED[3] ? 4 : (PL_LINK_CAP_MAX_LINK_SPEED[2] ? 3 : (PL_LINK_CAP_MAX_LINK_SPEED[1] ? 2 : 1))) ),                    
    .PHY_ASYNC_EN     ( ((PF0_LINK_STATUS_SLOT_CLOCK_CONFIG == "TRUE") ? "FALSE" : "TRUE" ) ),
    .PHY_REFCLK_FREQ  ( PHY_REFCLK_FREQ ),           
    .PHY_MCAPCLK_FREQ ( (((CRM_USER_CLK_FREQ == 2'b00) & (CRM_MCAP_CLK_FREQ == 1'b0)) ? 1 : 2) ),
    .PHY_USERCLK_FREQ ( (((CRM_USER_CLK_FREQ == 2'b10) | ((CRM_USER_CLK_FREQ == 2'b11) & (CRM_CORE_CLK_FREQ_500 == "TRUE"))) ? ((FPGA_XCVR == "HLF")? 2: 3) :
                                                                                                                               (CRM_USER_CLK_FREQ == 2'b01) ? 2 : 1) ),           
    .PHY_CORECLK_FREQ ( ((CRM_CORE_CLK_FREQ_500 == "TRUE") ? ((FPGA_XCVR == "HLF")? 1: 2) : 1) ) 
  ) gt_top_smsw_i (                                         

    //--------------------------------------------------------------------------
    //  Clock & Reset Ports
    //--------------------------------------------------------------------------
    .PHY_REFCLK          ( sys_clk_bufg ),      
    .PHY_USERCLK         ( user_clk ),  
    .PHY_MCAPCLK         ( mcap_clk ),  
    .PHY_GTREFCLK        ( sys_clk_gt ),               
    .PHY_RST_N           ( sys_rst_n ),           
   
    .PHY_PCLK            ( pipe_clk ),  
    .PHY_CORECLK         ( core_clk ), 
                            
                                               
    //--------------------------------------------------------------------------
    //  Serial Line Ports
    //--------------------------------------------------------------------------
    
    .PHY_RXP            ( pci_exp_rxp ),               
    .PHY_RXN            ( pci_exp_rxn ),               
                         
    .PHY_TXP            ( pci_exp_txp ),               
    .PHY_TXN            ( pci_exp_txn ),   
                                                                       
    //--------------------------------------------------------------------------
    //  TX Data Ports 
    //--------------------------------------------------------------------------
    
    .PHY_TXDATA         (PHY_TXDATA),            
    .PHY_TXDATAK        (PHY_TXDATAK),
    .PHY_TXDATA_VALID   (PHY_TXDATA_VALID),
    .PHY_TXSTART_BLOCK  (PHY_TXSTART_BLOCK),
    .PHY_TXSYNC_HEADER  (PHY_TXSYNC_HEADER), 

    //--------------------------------------------------------------------------
    //  RX Data Ports 
    //--------------------------------------------------------------------------

    .PHY_RXDATA         ( PHY_RXDATA ),
    .PHY_RXDATAK        ( PHY_RXDATAK ), 
    .PHY_RXDATA_VALID   ( PHY_RXDATA_VALID ),
    .PHY_RXSTART_BLOCK  ( PHY_RXSTART_BLOCK ), 
    .PHY_RXSYNC_HEADER  ( rxsync_header_nogate ),

    //--------------------------------------------------------------------------
    //  PHY Command Port
    //--------------------------------------------------------------------------
   
    .PHY_TXDETECTRX     ( pipe_tx_rcvr_det ),  
    .PHY_TXELECIDLE     (PHY_TXELECIDLE),                    
    .PHY_TXCOMPLIANCE   (PHY_TXCOMPLIANCE), 
    .PHY_RXPOLARITY     (PHY_RXPOLARITY),
    .PHY_POWERDOWN      ( pipe_tx00_powerdown ), 
    .PHY_RATE           ( pipe_tx_rate ),
    
    //--------------------------------------------------------------------------   
    //  PHY Status Ports
    //-------------------------------------------------------------------------- 
    
    .PHY_RXVALID        ( PHY_RXVALID  ),
    .PHY_PHYSTATUS      ( PHY_PHYSTATUS  ),
    .PHY_PHYSTATUS_RST  ( phy_rdy_phystatus ),
    .PHY_RXELECIDLE     ( PHY_RXELECIDLE ), 
    .PHY_RXSTATUS       ( PHY_RXSTATUS  ),
    
    //--------------------------------------------------------------------------
    //  TX Driver Ports
    //--------------------------------------------------------------------------
    
    .PHY_TXMARGIN       ( pipe_tx_margin ),          
    .PHY_TXSWING        ( pipe_tx_swing  ),           
    .PHY_TXDEEMPH       ( pipe_tx_deemph  ),    
    
    //--------------------------------------------------------------------------   
    //  TX Equalization Ports for Gen3
    //--------------------------------------------------------------------------  
    
    .PHY_TXEQ_CTRL      (PHY_TXEQ_CTRL),
    .PHY_TXEQ_PRESET    (PHY_TXEQ_PRESET),
    .PHY_TXEQ_COEFF     (PHY_TXEQ_COEFF), 
    .PHY_TXEQ_FS        ( pipe_eq_fs ),           
    .PHY_TXEQ_LF        ( pipe_eq_lf ),           
    .PHY_TXEQ_NEW_COEFF ( PHY_TXEQ_NEW_COEFF ),
    .PHY_TXEQ_DONE      ( PHY_TXEQ_DONE ),
                                                                 
    //--------------------------------------------------------------------------
    //  RX Equalization Ports for Gen3
    //--------------------------------------------------------------------------                                               
    
    .PHY_RXEQ_CTRL        (PHY_RXEQ_CTRL), 
    .PHY_RXEQ_TXPRESET    ( {PL_LINK_CAP_MAX_LINK_WIDTH{pipe_rx_eq_lp_tx_preset}} ),
    .PHY_RXEQ_PRESET_SEL  ( PHY_RXEQ_LFFS_SEL  ),
    .PHY_RXEQ_NEW_TXCOEFF ( PHY_RXEQ_NEW_TXCOEFF ),
    .PHY_RXEQ_DONE        ( PHY_RXEQ_DONE  ),
    .PHY_RXEQ_ADAPT_DONE  ( PHY_RXEQ_ADAPT_DONE ),

    //--------------------------------------------------------------------------
    //  Assist Signals
    //--------------------------------------------------------------------------

    .AS_MAC_IN_DETECT     ( as_mac_in_detect_ff1 ),
    .AS_CDR_HOLD_REQ      ( as_cdr_hold_req_ff1 )
);

 assign  common_commands_out = 17'd0;
 assign  pipe_tx_0_sigs = 70'd0; 
 assign  pipe_tx_1_sigs = 70'd0;
 assign  pipe_tx_2_sigs = 70'd0;
 assign  pipe_tx_3_sigs = 70'd0;
 assign  pipe_tx_4_sigs = 70'd0;
 assign  pipe_tx_5_sigs = 70'd0;
 assign  pipe_tx_6_sigs = 70'd0;
 assign  pipe_tx_7_sigs = 70'd0;
 assign  pipe_tx_8_sigs = 70'd0; 
 assign  pipe_tx_9_sigs = 70'd0;
 assign  pipe_tx_10_sigs = 70'd0;
 assign  pipe_tx_11_sigs = 70'd0;
 assign  pipe_tx_12_sigs = 70'd0;
 assign  pipe_tx_13_sigs = 70'd0;
 assign  pipe_tx_14_sigs = 70'd0;
 assign  pipe_tx_15_sigs = 70'd0;
 assign  phy_rdy = ~phy_rdy_phystatus;
end
endgenerate

assign { pipe_rx15_data[63:0], pipe_rx14_data[63:0], 
	       pipe_rx13_data[63:0], pipe_rx12_data[63:0],
	       pipe_rx11_data[63:0], pipe_rx10_data[63:0], 
	       pipe_rx09_data[63:0], pipe_rx08_data[63:0], 
	       pipe_rx07_data[63:0], pipe_rx06_data[63:0], 
	       pipe_rx05_data[63:0], pipe_rx04_data[63:0], 
         pipe_rx03_data[63:0], pipe_rx02_data[63:0], 
	       pipe_rx01_data[63:0], pipe_rx00_data[63:0]} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_RXDATA : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 64){1'b0}},PHY_RXDATA});

assign { pipe_rx15_char_is_k[1:0], pipe_rx14_char_is_k[1:0], 
	       pipe_rx13_char_is_k[1:0], pipe_rx12_char_is_k[1:0], 
         pipe_rx11_char_is_k[1:0], pipe_rx10_char_is_k[1:0], 
	       pipe_rx09_char_is_k[1:0], pipe_rx08_char_is_k[1:0], 
         pipe_rx07_char_is_k[1:0], pipe_rx06_char_is_k[1:0], 
	       pipe_rx05_char_is_k[1:0], pipe_rx04_char_is_k[1:0], 
         pipe_rx03_char_is_k[1:0], pipe_rx02_char_is_k[1:0], 
	       pipe_rx01_char_is_k[1:0], pipe_rx00_char_is_k[1:0]} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_RXDATAK : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 2){1'b0}},PHY_RXDATAK});

assign { pipe_rx15_data_valid, pipe_rx14_data_valid, 
	       pipe_rx13_data_valid, pipe_rx12_data_valid, 
         pipe_rx11_data_valid, pipe_rx10_data_valid, 
	       pipe_rx09_data_valid, pipe_rx08_data_valid, 
         pipe_rx07_data_valid, pipe_rx06_data_valid, 
	       pipe_rx05_data_valid, pipe_rx04_data_valid, 
         pipe_rx03_data_valid, pipe_rx02_data_valid, 
	       pipe_rx01_data_valid, pipe_rx00_data_valid} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_RXDATA_VALID : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 1){1'b0}},PHY_RXDATA_VALID});

assign { pipe_rx15_start_block[1:0], pipe_rx14_start_block[1:0], 
	       pipe_rx13_start_block[1:0], pipe_rx12_start_block[1:0], 
         pipe_rx11_start_block[1:0], pipe_rx10_start_block[1:0], 
	       pipe_rx09_start_block[1:0], pipe_rx08_start_block[1:0], 
         pipe_rx07_start_block[1:0], pipe_rx06_start_block[1:0], 
	       pipe_rx05_start_block[1:0], pipe_rx04_start_block[1:0], 
         pipe_rx03_start_block[1:0], pipe_rx02_start_block[1:0], 
	       pipe_rx01_start_block[1:0], pipe_rx00_start_block[1:0]} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_RXSTART_BLOCK : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 2){1'b0}},PHY_RXSTART_BLOCK});

assign { pipe_rx15_sync_header[1:0], pipe_rx14_sync_header[1:0], 
	       pipe_rx13_sync_header[1:0], pipe_rx12_sync_header[1:0], 
         pipe_rx11_sync_header[1:0], pipe_rx10_sync_header[1:0], 
	       pipe_rx09_sync_header[1:0], pipe_rx08_sync_header[1:0],
         pipe_rx07_sync_header[1:0], pipe_rx06_sync_header[1:0], 
	       pipe_rx05_sync_header[1:0], pipe_rx04_sync_header[1:0], 
         pipe_rx03_sync_header[1:0], pipe_rx02_sync_header[1:0], 
	       pipe_rx01_sync_header[1:0], pipe_rx00_sync_header[1:0]} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_RXSYNC_HEADER : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 2){1'b0}},PHY_RXSYNC_HEADER});

assign { pipe_rx15_valid, pipe_rx14_valid, 
	       pipe_rx13_valid, pipe_rx12_valid, 
         pipe_rx11_valid, pipe_rx10_valid, 
	       pipe_rx09_valid, pipe_rx08_valid, 
         pipe_rx07_valid, pipe_rx06_valid, 
	       pipe_rx05_valid, pipe_rx04_valid, 
         pipe_rx03_valid, pipe_rx02_valid, 
	       pipe_rx01_valid, pipe_rx00_valid} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_RXVALID : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 1){1'b0}},PHY_RXVALID});


// Soft fix to pass phystatus[0] (the last-done lane) to all other lanes in TO_2_DETECT state to make sure all other lanes are done.

always @(posedge pipe_clk or posedge sys_or_hot_rst) begin
   if (sys_or_hot_rst) begin
      pipe_tx_rate_ff   <= 2'b00;
   end else begin
      pipe_tx_rate_ff   <= pipe_tx_rate;
   end
end

always @(posedge pipe_clk or posedge sys_or_hot_rst) begin
   if (sys_or_hot_rst) begin
      speed_change_in_progress <= 1'b0;
   end else if (pipe_tx_rate != pipe_tx_rate_ff) begin
      speed_change_in_progress <= 1'b1;
   end else if (pipe_rx00_phy_status) begin
      speed_change_in_progress <= 1'b0;
   end
end

assign phy_status_fix   = (speed_change_in_progress)? {PL_LINK_CAP_MAX_LINK_WIDTH{PHY_PHYSTATUS[0]}}: PHY_PHYSTATUS;

assign { pipe_rx15_phy_status, pipe_rx14_phy_status, 
	       pipe_rx13_phy_status, pipe_rx12_phy_status, 
         pipe_rx11_phy_status, pipe_rx10_phy_status, 
	       pipe_rx09_phy_status, pipe_rx08_phy_status, 
         pipe_rx07_phy_status, pipe_rx06_phy_status, 
	       pipe_rx05_phy_status, pipe_rx04_phy_status, 
         pipe_rx03_phy_status, pipe_rx02_phy_status, 
	       pipe_rx01_phy_status, pipe_rx00_phy_status} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? phy_status_fix : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 1){1'b0}},phy_status_fix});

assign { pipe_rx15_elec_idle, pipe_rx14_elec_idle, pipe_rx13_elec_idle, pipe_rx12_elec_idle, 
         pipe_rx11_elec_idle, pipe_rx10_elec_idle, pipe_rx09_elec_idle, pipe_rx08_elec_idle, 
         pipe_rx07_elec_idle, pipe_rx06_elec_idle, pipe_rx05_elec_idle, pipe_rx04_elec_idle, 
         pipe_rx03_elec_idle, pipe_rx02_elec_idle, pipe_rx01_elec_idle, pipe_rx00_elec_idle} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_RXELECIDLE : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 1){1'b0}},PHY_RXELECIDLE});

assign { pipe_rx15_status, pipe_rx14_status, pipe_rx13_status, pipe_rx12_status, 
         pipe_rx11_status, pipe_rx10_status, pipe_rx09_status, pipe_rx08_status, 
         pipe_rx07_status, pipe_rx06_status, pipe_rx05_status, pipe_rx04_status, 
         pipe_rx03_status, pipe_rx02_status, pipe_rx01_status, pipe_rx00_status} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_RXSTATUS : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 3){1'b0}},PHY_RXSTATUS});

assign { pipe_tx15_eq_coeff, pipe_tx14_eq_coeff, 
	       pipe_tx13_eq_coeff, pipe_tx12_eq_coeff, 
         pipe_tx11_eq_coeff, pipe_tx10_eq_coeff, 
	       pipe_tx09_eq_coeff, pipe_tx08_eq_coeff, 
         pipe_tx07_eq_coeff, pipe_tx06_eq_coeff, 
	       pipe_tx05_eq_coeff, pipe_tx04_eq_coeff, 
         pipe_tx03_eq_coeff, pipe_tx02_eq_coeff, 
	       pipe_tx01_eq_coeff, pipe_tx00_eq_coeff} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_TXEQ_NEW_COEFF : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 18){1'b0}},PHY_TXEQ_NEW_COEFF});

assign { pipe_tx15_eq_done, pipe_tx14_eq_done, 
	       pipe_tx13_eq_done, pipe_tx12_eq_done, 
         pipe_tx11_eq_done, pipe_tx10_eq_done, 
	       pipe_tx09_eq_done, pipe_tx08_eq_done, 
         pipe_tx07_eq_done, pipe_tx06_eq_done, 
	       pipe_tx05_eq_done, pipe_tx04_eq_done, 
         pipe_tx03_eq_done, pipe_tx02_eq_done, 
	       pipe_tx01_eq_done, pipe_tx00_eq_done} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_TXEQ_DONE : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 1){1'b0}},PHY_TXEQ_DONE});

assign { pipe_rx15_eq_lp_lf_fs_sel, pipe_rx14_eq_lp_lf_fs_sel, 
	       pipe_rx13_eq_lp_lf_fs_sel, pipe_rx12_eq_lp_lf_fs_sel, 
         pipe_rx11_eq_lp_lf_fs_sel, pipe_rx10_eq_lp_lf_fs_sel, 
	       pipe_rx09_eq_lp_lf_fs_sel, pipe_rx08_eq_lp_lf_fs_sel, 
         pipe_rx07_eq_lp_lf_fs_sel, pipe_rx06_eq_lp_lf_fs_sel, 
	       pipe_rx05_eq_lp_lf_fs_sel, pipe_rx04_eq_lp_lf_fs_sel, 
         pipe_rx03_eq_lp_lf_fs_sel, pipe_rx02_eq_lp_lf_fs_sel, 
	       pipe_rx01_eq_lp_lf_fs_sel, pipe_rx00_eq_lp_lf_fs_sel} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_RXEQ_LFFS_SEL : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 1){1'b0}},PHY_RXEQ_LFFS_SEL});

assign { pipe_rx15_eq_lp_new_tx_coeff_or_preset, pipe_rx14_eq_lp_new_tx_coeff_or_preset, 
	       pipe_rx13_eq_lp_new_tx_coeff_or_preset, pipe_rx12_eq_lp_new_tx_coeff_or_preset, 
         pipe_rx11_eq_lp_new_tx_coeff_or_preset, pipe_rx10_eq_lp_new_tx_coeff_or_preset, 
	       pipe_rx09_eq_lp_new_tx_coeff_or_preset, pipe_rx08_eq_lp_new_tx_coeff_or_preset, 
         pipe_rx07_eq_lp_new_tx_coeff_or_preset, pipe_rx06_eq_lp_new_tx_coeff_or_preset, 
	       pipe_rx05_eq_lp_new_tx_coeff_or_preset, pipe_rx04_eq_lp_new_tx_coeff_or_preset, 
         pipe_rx03_eq_lp_new_tx_coeff_or_preset, pipe_rx02_eq_lp_new_tx_coeff_or_preset, 
	       pipe_rx01_eq_lp_new_tx_coeff_or_preset, pipe_rx00_eq_lp_new_tx_coeff_or_preset} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_RXEQ_NEW_TXCOEFF : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 18){1'b0}},PHY_RXEQ_NEW_TXCOEFF});

assign { pipe_rx15_eq_done, pipe_rx14_eq_done, pipe_rx13_eq_done, pipe_rx12_eq_done, 
         pipe_rx11_eq_done, pipe_rx10_eq_done, pipe_rx09_eq_done, pipe_rx08_eq_done, 
         pipe_rx07_eq_done, pipe_rx06_eq_done, pipe_rx05_eq_done, pipe_rx04_eq_done, 
         pipe_rx03_eq_done, pipe_rx02_eq_done, pipe_rx01_eq_done, pipe_rx00_eq_done} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_RXEQ_DONE : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 1){1'b0}},PHY_RXEQ_DONE});

assign { pipe_rx15_eq_lp_adapt_done, pipe_rx14_eq_lp_adapt_done, 
	       pipe_rx13_eq_lp_adapt_done, pipe_rx12_eq_lp_adapt_done, 
         pipe_rx11_eq_lp_adapt_done, pipe_rx10_eq_lp_adapt_done, 
	       pipe_rx09_eq_lp_adapt_done, pipe_rx08_eq_lp_adapt_done, 
         pipe_rx07_eq_lp_adapt_done, pipe_rx06_eq_lp_adapt_done, 
	       pipe_rx05_eq_lp_adapt_done, pipe_rx04_eq_lp_adapt_done, 
         pipe_rx03_eq_lp_adapt_done, pipe_rx02_eq_lp_adapt_done, 
	       pipe_rx01_eq_lp_adapt_done, pipe_rx00_eq_lp_adapt_done} = (PL_LINK_CAP_MAX_LINK_WIDTH == 16 ? PHY_RXEQ_ADAPT_DONE : {{((16-PL_LINK_CAP_MAX_LINK_WIDTH) * 1){1'b0}},PHY_RXEQ_ADAPT_DONE});

assign   sys_rst_n = sys_reset; //pcie_perst0_b; // Use the reset from pcie_4_0_pipe
assign   mcap_rst_b = ~sys_reset;
assign   user_lnk_up_int = (cfg_phy_link_status == 2'b11) ? 1'b1 : 1'b0;
assign   sys_or_hot_rst = ~sys_rst_n || cfg_hot_reset_out;

always @(posedge user_clk) begin

  if (!sys_rst_n) begin

    reg_user_lnk_up <= #TCQ 1'b0;

  end else begin

    reg_user_lnk_up <= #TCQ user_lnk_up_int;

  end

end
assign     user_lnk_up = reg_user_lnk_up;

always @(posedge user_clk or posedge sys_or_hot_rst) begin

  if (sys_or_hot_rst) begin

    user_reset_int <= #TCQ 1'b1;

  end else if (cfg_phy_link_status[1] && !cfg_phy_link_down) begin

    user_reset_int <= #TCQ 1'b0;
    
   end else if (cfg_phy_link_down) begin

    user_reset_int <= #TCQ 1'b1;
  end

end

always @(posedge user_clk or posedge sys_or_hot_rst) begin

  if (sys_or_hot_rst) begin

    reg_user_reset <= #TCQ 1'b1;

  end else begin

    reg_user_reset <= #TCQ user_reset_int;

  end

end
assign user_reset = reg_user_reset;


assign PHY_TXDATA = ( PL_LINK_CAP_MAX_LINK_WIDTH==16 ?
                         { 32'h0, pipe_tx15_data[31:0], 32'h0, pipe_tx14_data[31:0], 
			                     32'h0, pipe_tx13_data[31:0], 32'h0, pipe_tx12_data[31:0], 
			                     32'h0, pipe_tx11_data[31:0], 32'h0, pipe_tx10_data[31:0], 
			                     32'h0, pipe_tx09_data[31:0], 32'h0, pipe_tx08_data[31:0], 
			                     pipe_tx15_data[31:0], pipe_tx07_data[31:0], pipe_tx14_data[31:0], pipe_tx06_data[31:0],
                           pipe_tx13_data[31:0], pipe_tx05_data[31:0], pipe_tx12_data[31:0], pipe_tx04_data[31:0], 
                           pipe_tx11_data[31:0], pipe_tx03_data[31:0], pipe_tx10_data[31:0], pipe_tx02_data[31:0],
                           pipe_tx09_data[31:0], pipe_tx01_data[31:0], pipe_tx08_data[31:0], pipe_tx00_data[31:0]} :
                      PL_LINK_CAP_MAX_LINK_WIDTH==8 ?
			                   { pipe_tx15_data[31:0], pipe_tx07_data[31:0], pipe_tx14_data[31:0], pipe_tx06_data[31:0], 
			                     pipe_tx13_data[31:0], pipe_tx05_data[31:0], pipe_tx12_data[31:0], pipe_tx04_data[31:0], 
                           pipe_tx11_data[31:0], pipe_tx03_data[31:0], pipe_tx10_data[31:0], pipe_tx02_data[31:0], 
			                     pipe_tx09_data[31:0], pipe_tx01_data[31:0], pipe_tx08_data[31:0], pipe_tx00_data[31:0]} :
                      PL_LINK_CAP_MAX_LINK_WIDTH==4 ?
			                   { pipe_tx11_data[31:0], pipe_tx03_data[31:0], pipe_tx10_data[31:0], pipe_tx02_data[31:0], 
			                     pipe_tx09_data[31:0], pipe_tx01_data[31:0], pipe_tx08_data[31:0], pipe_tx00_data[31:0]} :
                      PL_LINK_CAP_MAX_LINK_WIDTH==2 ?
			                   { pipe_tx09_data[31:0], pipe_tx01_data[31:0], pipe_tx08_data[31:0], pipe_tx00_data[31:0]} : 
			                   {pipe_tx08_data[31:0], pipe_tx00_data[31:0]} );            

 assign PHY_TXDATAK = ( PL_LINK_CAP_MAX_LINK_WIDTH==16 ?
                         { pipe_tx15_char_is_k[1:0], pipe_tx14_char_is_k[1:0], pipe_tx13_char_is_k[1:0], pipe_tx12_char_is_k[1:0], 
                           pipe_tx11_char_is_k[1:0], pipe_tx10_char_is_k[1:0], pipe_tx09_char_is_k[1:0], pipe_tx08_char_is_k[1:0], 
                           pipe_tx07_char_is_k[1:0], pipe_tx06_char_is_k[1:0], pipe_tx05_char_is_k[1:0], pipe_tx04_char_is_k[1:0], 
                           pipe_tx03_char_is_k[1:0], pipe_tx02_char_is_k[1:0], pipe_tx01_char_is_k[1:0], pipe_tx00_char_is_k[1:0]} :
                        PL_LINK_CAP_MAX_LINK_WIDTH==8 ?
                         { pipe_tx07_char_is_k[1:0], pipe_tx06_char_is_k[1:0], pipe_tx05_char_is_k[1:0], pipe_tx04_char_is_k[1:0], 
                           pipe_tx03_char_is_k[1:0], pipe_tx02_char_is_k[1:0], pipe_tx01_char_is_k[1:0], pipe_tx00_char_is_k[1:0]} :
                        PL_LINK_CAP_MAX_LINK_WIDTH==4 ?
                         { pipe_tx03_char_is_k[1:0], pipe_tx02_char_is_k[1:0], pipe_tx01_char_is_k[1:0], pipe_tx00_char_is_k[1:0]} :
                        PL_LINK_CAP_MAX_LINK_WIDTH==2 ?
                         { pipe_tx01_char_is_k[1:0], pipe_tx00_char_is_k[1:0]} : pipe_tx00_char_is_k[1:0] );

assign PHY_TXDATA_VALID = ( PL_LINK_CAP_MAX_LINK_WIDTH==16 ?
                         { pipe_tx15_data_valid, pipe_tx14_data_valid, pipe_tx13_data_valid, pipe_tx12_data_valid, 
                           pipe_tx11_data_valid, pipe_tx10_data_valid, pipe_tx09_data_valid, pipe_tx08_data_valid, 
                           pipe_tx07_data_valid, pipe_tx06_data_valid, pipe_tx05_data_valid, pipe_tx04_data_valid, 
                           pipe_tx03_data_valid, pipe_tx02_data_valid, pipe_tx01_data_valid, pipe_tx00_data_valid} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==8 ?
                         { pipe_tx07_data_valid, pipe_tx06_data_valid, pipe_tx05_data_valid, pipe_tx04_data_valid, 
                           pipe_tx03_data_valid, pipe_tx02_data_valid, pipe_tx01_data_valid, pipe_tx00_data_valid} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==4 ?
                         { pipe_tx03_data_valid, pipe_tx02_data_valid, pipe_tx01_data_valid, pipe_tx00_data_valid} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==2 ?
                         { pipe_tx01_data_valid, pipe_tx00_data_valid} : pipe_tx00_data_valid );

assign PHY_TXSTART_BLOCK = ( PL_LINK_CAP_MAX_LINK_WIDTH==16 ?
                         { pipe_tx15_start_block, pipe_tx15_start_block, pipe_tx15_start_block, pipe_tx15_start_block, 
                           pipe_tx11_start_block, pipe_tx10_start_block, pipe_tx09_start_block, pipe_tx08_start_block,                      
                           pipe_tx07_start_block, pipe_tx06_start_block, pipe_tx05_start_block, pipe_tx04_start_block, 
                           pipe_tx03_start_block, pipe_tx02_start_block, pipe_tx01_start_block, pipe_tx00_start_block} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==8 ?
                         { pipe_tx07_start_block, pipe_tx06_start_block, pipe_tx05_start_block, pipe_tx04_start_block, 
                           pipe_tx03_start_block, pipe_tx02_start_block, pipe_tx01_start_block, pipe_tx00_start_block} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==4 ?
                         { pipe_tx03_start_block, pipe_tx02_start_block, pipe_tx01_start_block, pipe_tx00_start_block} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==2 ?
                         { pipe_tx01_start_block, pipe_tx00_start_block} : pipe_tx00_start_block );

assign PHY_TXSYNC_HEADER = ( PL_LINK_CAP_MAX_LINK_WIDTH==16 ?
                         { pipe_tx15_sync_header[1:0], pipe_tx14_sync_header[1:0], pipe_tx13_sync_header[1:0], pipe_tx12_sync_header[1:0], 
                           pipe_tx11_sync_header[1:0], pipe_tx10_sync_header[1:0], pipe_tx09_sync_header[1:0], pipe_tx08_sync_header[1:0],
                           pipe_tx07_sync_header[1:0], pipe_tx06_sync_header[1:0], pipe_tx05_sync_header[1:0], pipe_tx04_sync_header[1:0], 
                           pipe_tx03_sync_header[1:0], pipe_tx02_sync_header[1:0], pipe_tx01_sync_header[1:0], pipe_tx00_sync_header[1:0]} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==8 ?
                         { pipe_tx07_sync_header[1:0], pipe_tx06_sync_header[1:0], pipe_tx05_sync_header[1:0], pipe_tx04_sync_header[1:0], 
                           pipe_tx03_sync_header[1:0], pipe_tx02_sync_header[1:0], pipe_tx01_sync_header[1:0], pipe_tx00_sync_header[1:0]} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==4 ?
                         { pipe_tx03_sync_header[1:0], pipe_tx02_sync_header[1:0], pipe_tx01_sync_header[1:0], pipe_tx00_sync_header[1:0]} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==2 ?
                         { pipe_tx01_sync_header[1:0], pipe_tx00_sync_header[1:0]} : pipe_tx00_sync_header[1:0] );

assign PHY_TXELECIDLE = ( PL_LINK_CAP_MAX_LINK_WIDTH==16 ?
                        { pipe_tx15_elec_idle, pipe_tx14_elec_idle, pipe_tx13_elec_idle, pipe_tx12_elec_idle, 
                          pipe_tx11_elec_idle, pipe_tx10_elec_idle, pipe_tx09_elec_idle, pipe_tx08_elec_idle, 
                          pipe_tx07_elec_idle, pipe_tx06_elec_idle, pipe_tx05_elec_idle, pipe_tx04_elec_idle, 
                          pipe_tx03_elec_idle, pipe_tx02_elec_idle, pipe_tx01_elec_idle, pipe_tx00_elec_idle} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==8 ?
                        { pipe_tx07_elec_idle, pipe_tx06_elec_idle, pipe_tx05_elec_idle, pipe_tx04_elec_idle, 
                          pipe_tx03_elec_idle, pipe_tx02_elec_idle, pipe_tx01_elec_idle, pipe_tx00_elec_idle} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==4 ?
                        { pipe_tx03_elec_idle, pipe_tx02_elec_idle, pipe_tx01_elec_idle, pipe_tx00_elec_idle} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==2 ?
                        { pipe_tx01_elec_idle, pipe_tx00_elec_idle} : pipe_tx00_elec_idle );


assign PHY_TXCOMPLIANCE = ( PL_LINK_CAP_MAX_LINK_WIDTH==16 ?
                        { pipe_tx15_compliance, pipe_tx14_compliance, pipe_tx13_compliance, pipe_tx12_compliance, 
                          pipe_tx11_compliance, pipe_tx10_compliance, pipe_tx09_compliance, pipe_tx08_compliance, 
                          pipe_tx07_compliance, pipe_tx06_compliance, pipe_tx05_compliance, pipe_tx04_compliance, 
                          pipe_tx03_compliance, pipe_tx02_compliance, pipe_tx01_compliance, pipe_tx00_compliance} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==8 ?
                        { pipe_tx07_compliance, pipe_tx06_compliance, pipe_tx05_compliance, pipe_tx04_compliance, 
                          pipe_tx03_compliance, pipe_tx02_compliance, pipe_tx01_compliance, pipe_tx00_compliance} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==4 ?
                        { pipe_tx03_compliance, pipe_tx02_compliance, pipe_tx01_compliance, pipe_tx00_compliance} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==2 ?
                        { pipe_tx01_compliance, pipe_tx00_compliance} : pipe_tx00_compliance );

assign PHY_RXPOLARITY =  ( 
                          PL_LINK_CAP_MAX_LINK_WIDTH==16 ?
                        { pipe_rx15_polarity, pipe_rx14_polarity, pipe_rx13_polarity, pipe_rx12_polarity, 
                          pipe_rx11_polarity, pipe_rx10_polarity, pipe_rx09_polarity, pipe_rx08_polarity, 
                          pipe_rx07_polarity, pipe_rx06_polarity, pipe_rx05_polarity, pipe_rx04_polarity, 
                          pipe_rx03_polarity, pipe_rx02_polarity, pipe_rx01_polarity, pipe_rx00_polarity} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==8 ?
                        { pipe_rx07_polarity, pipe_rx06_polarity, pipe_rx05_polarity, pipe_rx04_polarity, 
                          pipe_rx03_polarity, pipe_rx02_polarity, pipe_rx01_polarity, pipe_rx00_polarity} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==4 ?
                        { pipe_rx03_polarity, pipe_rx02_polarity, pipe_rx01_polarity, pipe_rx00_polarity} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==2 ?
                        { pipe_rx01_polarity, pipe_rx00_polarity} : pipe_rx00_polarity );

assign PHY_TXEQ_CTRL = ( PL_LINK_CAP_MAX_LINK_WIDTH==16 ? 
                          { pipe_tx15_eq_control, pipe_tx14_eq_control, pipe_tx13_eq_control, pipe_tx12_eq_control, 
			    pipe_tx11_eq_control, pipe_tx10_eq_control, pipe_tx09_eq_control, pipe_tx08_eq_control, 
			    pipe_tx07_eq_control, pipe_tx06_eq_control, pipe_tx05_eq_control, pipe_tx04_eq_control, 
                            pipe_tx03_eq_control, pipe_tx02_eq_control, pipe_tx01_eq_control, pipe_tx00_eq_control} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==8 ?
                          { pipe_tx07_eq_control, pipe_tx06_eq_control, pipe_tx05_eq_control, pipe_tx04_eq_control, 
                            pipe_tx03_eq_control, pipe_tx02_eq_control, pipe_tx01_eq_control, pipe_tx00_eq_control} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==4 ?
                          { pipe_tx03_eq_control, pipe_tx02_eq_control, pipe_tx01_eq_control, pipe_tx00_eq_control} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==2 ?
                          { pipe_tx01_eq_control, pipe_tx00_eq_control} : pipe_tx00_eq_control );

assign PHY_TXEQ_PRESET = (  PL_LINK_CAP_MAX_LINK_WIDTH==16 ?
                          { pipe_tx15_eq_deemph[3:0], pipe_tx14_eq_deemph[3:0], pipe_tx13_eq_deemph[3:0], pipe_tx12_eq_deemph[3:0],
                            pipe_tx11_eq_deemph[3:0], pipe_tx10_eq_deemph[3:0], pipe_tx09_eq_deemph[3:0], pipe_tx08_eq_deemph[3:0],
                            pipe_tx07_eq_deemph[3:0], pipe_tx06_eq_deemph[3:0], pipe_tx05_eq_deemph[3:0], pipe_tx04_eq_deemph[3:0],
                            pipe_tx03_eq_deemph[3:0], pipe_tx02_eq_deemph[3:0], pipe_tx01_eq_deemph[3:0], pipe_tx00_eq_deemph[3:0]} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==8 ?
                          { pipe_tx07_eq_deemph[3:0], pipe_tx06_eq_deemph[3:0], pipe_tx05_eq_deemph[3:0], pipe_tx04_eq_deemph[3:0],
                            pipe_tx03_eq_deemph[3:0], pipe_tx02_eq_deemph[3:0], pipe_tx01_eq_deemph[3:0], pipe_tx00_eq_deemph[3:0]} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==4 ?
                          { pipe_tx03_eq_deemph[3:0], pipe_tx02_eq_deemph[3:0], pipe_tx01_eq_deemph[3:0], pipe_tx00_eq_deemph[3:0]} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==2 ?
                          { pipe_tx01_eq_deemph[3:0], pipe_tx00_eq_deemph[3:0]} :  pipe_tx00_eq_deemph[3:0] );

assign PHY_TXEQ_COEFF = ( PL_LINK_CAP_MAX_LINK_WIDTH==16 ?
                          { pipe_tx15_eq_deemph, pipe_tx14_eq_deemph, pipe_tx13_eq_deemph, pipe_tx12_eq_deemph,
                            pipe_tx11_eq_deemph, pipe_tx10_eq_deemph, pipe_tx09_eq_deemph, pipe_tx08_eq_deemph,
                            pipe_tx07_eq_deemph, pipe_tx06_eq_deemph, pipe_tx05_eq_deemph, pipe_tx04_eq_deemph,
                            pipe_tx03_eq_deemph, pipe_tx02_eq_deemph, pipe_tx01_eq_deemph, pipe_tx00_eq_deemph} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==8 ?
                          { pipe_tx07_eq_deemph, pipe_tx06_eq_deemph, pipe_tx05_eq_deemph, pipe_tx04_eq_deemph,
                            pipe_tx03_eq_deemph, pipe_tx02_eq_deemph, pipe_tx01_eq_deemph, pipe_tx00_eq_deemph} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==4 ?
                          { pipe_tx03_eq_deemph, pipe_tx02_eq_deemph, pipe_tx01_eq_deemph, pipe_tx00_eq_deemph} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==2 ?
                          { pipe_tx01_eq_deemph, pipe_tx00_eq_deemph} : pipe_tx00_eq_deemph );

assign PHY_RXEQ_CTRL = ( PL_LINK_CAP_MAX_LINK_WIDTH==16 ?
                          { pipe_rx15_eq_control, pipe_rx14_eq_control, pipe_rx13_eq_control, pipe_rx12_eq_control, 
                            pipe_rx11_eq_control, pipe_rx10_eq_control, pipe_rx09_eq_control, pipe_rx08_eq_control, 
                            pipe_rx07_eq_control, pipe_rx06_eq_control, pipe_rx05_eq_control, pipe_rx04_eq_control, 
                            pipe_rx03_eq_control, pipe_rx02_eq_control, pipe_rx01_eq_control, pipe_rx00_eq_control} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==8 ?
                          { pipe_rx07_eq_control, pipe_rx06_eq_control, pipe_rx05_eq_control, pipe_rx04_eq_control, 
                            pipe_rx03_eq_control, pipe_rx02_eq_control, pipe_rx01_eq_control, pipe_rx00_eq_control} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==4 ?
                          { pipe_rx03_eq_control, pipe_rx02_eq_control, pipe_rx01_eq_control, pipe_rx00_eq_control} :
                          PL_LINK_CAP_MAX_LINK_WIDTH==2 ?
                          { pipe_rx01_eq_control, pipe_rx00_eq_control} : pipe_rx00_eq_control );

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_phy_top.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
/*****************************************************************************
** Description:
**    PCIe Gen4 PHY supports:
**       - Gen1: per-lane 16b @ 125MHz
**       - Gen2: per-lane 16b @ 250MHz
**       - Gen3: per-lane 32b @ 250Mhz
**       - Gen4: per-lane 64b @ 250MHz
**
******************************************************************************/
//--------------------------------------------------------------------------------------------------
//  Design :  PHY Wrapper
//  Module :  PHY Wrapper
//--------------------------------------------------------------------------------------------------

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_phy_top #(
   // Parameters
   parameter         FPGA_FAMILY       = "US",     // "US" = UltraScale; "USM" = Diablo
   parameter         FPGA_XCVR         = "H",      // "H" = GTH; "Y" = GTY; "Y64" = GTY-64b
   parameter integer PIPELINE_STAGES   = 0,        // 0 = no pipeline; 1 = 1 stage; 2 = 2 stages; 3 = 3 stages
   parameter         PHY_SIM_EN        = "FALSE",  // "FALSE" = Normal; "TRUE"  = Simulation
   parameter integer PHY_LANE          = 1,        // Valid settings: 1, 2, 4, 8, 16(only for Gen1/2/3)
   parameter integer PHY_MAX_SPEED     = 3,        // 1 = Gen1 Capable; 2 = Gen2 Capable; 3 = Gen3 Capable; 4 = Gen4 Capable   
   parameter         PHY_ASYNC_EN      = "FALSE",  // "FALSE" = Sync Clocking; "TRUE"  = Async Clocking
   parameter         PHY_REFCLK_FREQ   = 0,        // 0 = 100 MHz; 1 = 125 MHz; 2 = 250 MHz
   parameter integer PHY_CORECLK_FREQ  = 2,        // 1 = 250 MHz; 2 = 500 MHz
   parameter integer PHY_USERCLK_FREQ  = 3,        // 1 = 62.5 MHz; 2 = 125 MHz; 3 = 250 MHz; 4 = 500 MHz
   parameter integer PHY_MCAPCLK_FREQ  = 2,        // 1 = 62.5 MHz; 2 = 125 MHz
   parameter integer PHY_GT_TXPRESET   = 0,        // Valid settings: 0 to 10
   parameter integer PHY_LP_TXPRESET   = 5         // Valid settings: 5
)  (                                                         
   // Clock & Reset
   input  wire                         PHY_REFCLK,          
   input  wire                         PHY_GTREFCLK,     
   input  wire                         PHY_RST_N,           
   
   output wire                         PHY_CORECLK, 
   output wire                         PHY_USERCLK,                          
   output wire                         PHY_MCAPCLK,                          
   output wire                         PHY_PCLK,  
  
   // TX Data 
   input  wire [(PHY_LANE*64)-1:0]     PHY_TXDATA,            
   input  wire [(PHY_LANE* 2)-1:0]     PHY_TXDATAK,    
   input  wire [PHY_LANE-1:0]          PHY_TXDATA_VALID,
   input  wire [PHY_LANE-1:0]          PHY_TXSTART_BLOCK,      
   input  wire [(PHY_LANE* 2)-1:0]     PHY_TXSYNC_HEADER,                    

   output wire [PHY_LANE-1:0]          PHY_TXP,    // Serial Line      
   output wire [PHY_LANE-1:0]          PHY_TXN,    // Serial Line  

   // RX Data
   input  wire [PHY_LANE-1:0]          PHY_RXP,    // Serial Line           
   input  wire [PHY_LANE-1:0]          PHY_RXN,    // Serial Line

   output wire [(PHY_LANE*64)-1:0]     PHY_RXDATA,            
   output wire [(PHY_LANE* 2)-1:0]     PHY_RXDATAK,       
   output wire [PHY_LANE-1:0]          PHY_RXDATA_VALID,         
   output wire [(PHY_LANE* 2)-1:0]     PHY_RXSTART_BLOCK,        
   output wire [(PHY_LANE* 2)-1:0]     PHY_RXSYNC_HEADER,        

   // PHY Command
   input  wire                         PHY_TXDETECTRX,        
   input  wire [PHY_LANE-1:0]          PHY_TXELECIDLE,        
   input  wire [PHY_LANE-1:0]          PHY_TXCOMPLIANCE,      
   input  wire [PHY_LANE-1:0]          PHY_RXPOLARITY,        
   input  wire [1:0]                   PHY_POWERDOWN,         
   input  wire [1:0]                   PHY_RATE,              
    
   // PHY Status
   output wire [PHY_LANE-1:0]          PHY_RXVALID,               
   output wire [PHY_LANE-1:0]          PHY_PHYSTATUS,          
   output wire                         PHY_PHYSTATUS_RST,         
   output wire [PHY_LANE-1:0]          PHY_RXELECIDLE,         
   output wire [(PHY_LANE*3)-1:0]      PHY_RXSTATUS,                       
    
   // TX Driver
   input  wire [ 2:0]                  PHY_TXMARGIN,          
   input  wire                         PHY_TXSWING,           
   input  wire                         PHY_TXDEEMPH,    
    
   // TX Equalization (Gen3/4)
   input  wire [(PHY_LANE*2)-1:0]      PHY_TXEQ_CTRL,      
   input  wire [(PHY_LANE*4)-1:0]      PHY_TXEQ_PRESET,       
   input  wire [(PHY_LANE*6)-1:0]      PHY_TXEQ_COEFF,                                                            

   output wire [ 5:0]                  PHY_TXEQ_FS,           
   output wire [ 5:0]                  PHY_TXEQ_LF,           
   output wire [(PHY_LANE*18)-1:0]     PHY_TXEQ_NEW_COEFF,        
   output wire [PHY_LANE-1:0]          PHY_TXEQ_DONE,         

   // RX Equalization (Gen3/4)
   input  wire [(PHY_LANE*2)-1:0]      PHY_RXEQ_CTRL,     
   input  wire [(PHY_LANE*4)-1:0]      PHY_RXEQ_TXPRESET,      

   output wire [PHY_LANE-1:0]          PHY_RXEQ_PRESET_SEL,    
   output wire [(PHY_LANE*18)-1:0]     PHY_RXEQ_NEW_TXCOEFF,   
   output wire [PHY_LANE-1:0]          PHY_RXEQ_ADAPT_DONE,     
   output wire [PHY_LANE-1:0]          PHY_RXEQ_DONE,

   // Assist Signals
   input  wire                         AS_MAC_IN_DETECT,
   input  wire                         AS_CDR_HOLD_REQ
   );

   localparam  TCQ   = 1;

   wire                 phy_userclk_int;
   wire                 phy_mcapclk_int;
   wire                 phy_pclk;
   wire                 phy_pclk2;
   wire  [PHY_LANE-1:0]          phy_rxvalid_pclk2;
   wire  [PHY_LANE-1:0]          phy_phystatus_pclk2;
   wire                 phy_phystatus_rst_pclk2;
   wire  [(PHY_LANE* 3)-1:0]     phy_rxstatus_pclk2;
   wire  [5:0]          phy_txeq_fs_pclk2;
   wire  [5:0]          phy_txeq_lf_pclk2;
   wire  [(PHY_LANE* 18)-1:0]    phy_txeq_new_coeff_pclk2;
   wire  [PHY_LANE-1:0]          phy_txeq_done_pclk2;
   wire  [PHY_LANE-1:0]          phy_rxeq_preset_sel_pclk2;
   wire  [(PHY_LANE* 18)-1:0]    phy_rxeq_new_txcoeff_pclk2;
   wire  [PHY_LANE-1:0]          phy_rxeq_done_pclk2;
   wire  [PHY_LANE-1:0]          phy_rxeq_adapt_done_pclk2;

   wire                 phy_txdetectrx_32b;
   wire  [PHY_LANE-1:0]          phy_txelecidle_32b;
   wire  [PHY_LANE-1:0]          phy_txcompliance_32b;
   wire  [PHY_LANE-1:0]          phy_rxpolarity_32b;
   wire  [1:0]          phy_powerdown_32b;
   wire  [1:0]          phy_rate_32b;

   wire  [(PHY_LANE*32)-1:0]     phy_txdata_32b;            
   wire  [(PHY_LANE* 2)-1:0]     phy_txdatak_32b;            
   wire  [PHY_LANE-1:0]          phy_txdata_valid_32b;
   wire  [PHY_LANE-1:0]          phy_txstart_block_32b;      
   wire  [(PHY_LANE* 2)-1:0]     phy_txsync_header_32b;  
   wire  [(PHY_LANE*2)-1:0]      phy_txeq_ctrl_pclk2;            
   wire  [(PHY_LANE*4)-1:0]      phy_txeq_preset_pclk2;            
   wire  [(PHY_LANE*6)-1:0]      phy_txeq_coeff_pclk2;

   wire  [(PHY_LANE*64)-1:0]     phy_txdata_64b;            

   wire  [(PHY_LANE*32)-1:0]     phy_rxdata_32b;            
   wire  [(PHY_LANE* 2)-1:0]     phy_rxdatak_32b;            
   wire  [PHY_LANE-1:0]          phy_rxdata_valid_32b;
   wire  [PHY_LANE-1:0]          phy_rxstart_block_32b;      
   wire  [(PHY_LANE* 2)-1:0]     phy_rxsync_header_32b; 

   wire  [(PHY_LANE*64)-1:0]     phy_rxdata_64b;            
   wire  [(PHY_LANE* 2)-1:0]     phy_rxstart_block_64b;      

   wire  [(PHY_LANE*64)-1:0]     phy_txdata_pl;            
   wire  [(PHY_LANE* 2)-1:0]     phy_txdatak_pl;            
   wire  [PHY_LANE-1:0]          phy_txdata_valid_pl;
   wire  [PHY_LANE-1:0]          phy_txstart_block_pl;      
   wire  [(PHY_LANE* 2)-1:0]     phy_txsync_header_pl;  

   wire  [(PHY_LANE*64)-1:0]     phy_rxdata_pl;            
   wire  [(PHY_LANE* 2)-1:0]     phy_rxdatak_pl;            
   wire  [PHY_LANE-1:0]          phy_rxdata_valid_pl;
   wire  [(PHY_LANE* 2)-1:0]     phy_rxstart_block_pl;      
   wire  [(PHY_LANE* 2)-1:0]     phy_rxsync_header_pl; 

   wire                 phy_txdetectrx_pl;        
   wire  [PHY_LANE-1:0]          phy_txelecidle_pl;        
   wire  [PHY_LANE-1:0]          phy_txcompliance_pl;      
   wire  [PHY_LANE-1:0]          phy_rxpolarity_pl;        
   wire  [1:0]          phy_powerdown_pl;         
   wire  [1:0]          phy_rate_pl;   

   wire  [PHY_LANE-1:0]          phy_rxvalid_pl;               
   wire  [PHY_LANE-1:0]          phy_phystatus_pl;          
   wire  [PHY_LANE-1:0]          phy_rxelecidle_pl;         
   wire  [(PHY_LANE*3)-1:0]      phy_rxstatus_pl;          

   wire  [ 2:0]         phy_txmargin_pl;          
   wire                 phy_txswing_pl;           
   wire                 phy_txdeemph_pl;  

   wire  [(PHY_LANE*2)-1:0]      phy_txeq_ctrl_pl;      
   wire  [(PHY_LANE*4)-1:0]      phy_txeq_preset_pl;       
   wire  [(PHY_LANE*6)-1:0]      phy_txeq_coeff_pl;                                                            

   wire  [ 5:0]         phy_txeq_fs_pl;           
   wire  [ 5:0]         phy_txeq_lf_pl;           
   wire  [(PHY_LANE*18)-1:0]     phy_txeq_new_coeff_pl;        
   wire  [PHY_LANE-1:0]          phy_txeq_done_pl;         

   wire  [(PHY_LANE*2)-1:0]      phy_rxeq_ctrl_pl;     
   wire  [(PHY_LANE*4)-1:0]      phy_rxeq_txpreset_pl;      

   wire  [PHY_LANE-1:0]          phy_rxeq_preset_sel_pl;    
   wire  [(PHY_LANE*18)-1:0]     phy_rxeq_new_txcoeff_pl;   
   wire  [PHY_LANE-1:0]          phy_rxeq_adapt_done_pl;     
   wire  [PHY_LANE-1:0]          phy_rxeq_done_pl;

   wire                 as_mac_in_detect_pl;
   wire                 as_cdr_hold_req_pl;

   wire  [PHY_LANE-1:0]          com_det_lower;
   wire  [PHY_LANE-1:0]          com_det_upper;
   wire  [PHY_LANE-1:0]          idl_det_lower;
   wire  [PHY_LANE-1:0]          idl_det_upper;
   wire  [PHY_LANE-1:0]          eios_det_c0;
   wire  [PHY_LANE-1:0]          eios_det_c1;
   wire  [PHY_LANE-1:0]          eios_det_c2;
   wire  [PHY_LANE-1:0]          eios_det_c3;
   wire  [(PHY_LANE* 3)-1:0]     phy_rxstatus_raw;

   reg                  phy_rxelecidle_ff;
   reg                  phy_rxelecidle_ff2;
   reg                  phy_rxcdrhold_wire;
   reg                  phy_rxcdrhold_pclk2;

   reg   [PHY_LANE-1:0]          phy_rxstatus_mask_wire, phy_rxstatus_mask;
   reg   [PHY_LANE-1:0]          saved_com_det_lower_wire, saved_com_det_lower;
   reg   [PHY_LANE-1:0]          saved_com_det_upper_wire, saved_com_det_upper;

   //--------------------------------------------------------------------------
   //  Pipeline Stages
   //--------------------------------------------------------------------------        
   (* keep = "true", max_fanout = 500 *) wire   phy_phystatus_rst_int;
   assign phy_phystatus_rst_int  = PHY_PHYSTATUS_RST;

      // Programmable stages to ease GT lane routing
      xp4_usp_smsw_phy_pipeline #(
         //  Parameters
         .PIPELINE_STAGES  ( PIPELINE_STAGES ),
         .PHY_LANE         ( PHY_LANE ),
         .TCQ              ( TCQ )
      ) phy_pipeline_smsw (                                         
         // Clock & Reset Ports
         .phy_pclk               ( PHY_PCLK ),  
         .phy_rst                ( phy_phystatus_rst_int ),  

         // TX Data
         .phy_txdata_i           ( PHY_TXDATA ),
         .phy_txdatak_i          ( PHY_TXDATAK ),
         .phy_txdata_valid_i     ( PHY_TXDATA_VALID ),
         .phy_txstart_block_i    ( PHY_TXSTART_BLOCK ),
         .phy_txsync_header_i    ( PHY_TXSYNC_HEADER ),

         .phy_txdata_o           ( phy_txdata_pl ),
         .phy_txdatak_o          ( phy_txdatak_pl ),
         .phy_txdata_valid_o     ( phy_txdata_valid_pl ),
         .phy_txstart_block_o    ( phy_txstart_block_pl ),
         .phy_txsync_header_o    ( phy_txsync_header_pl ),

         // RX Data
         .phy_rxdata_i           ( phy_rxdata_pl ),            
         .phy_rxdatak_i          ( phy_rxdatak_pl ),       
         .phy_rxdata_valid_i     ( phy_rxdata_valid_pl ),         
         .phy_rxstart_block_i    ( phy_rxstart_block_pl ),        
         .phy_rxsync_header_i    ( phy_rxsync_header_pl ),   

         .phy_rxdata_o           ( PHY_RXDATA ),            
         .phy_rxdatak_o          ( PHY_RXDATAK ),       
         .phy_rxdata_valid_o     ( PHY_RXDATA_VALID ),         
         .phy_rxstart_block_o    ( PHY_RXSTART_BLOCK ),        
         .phy_rxsync_header_o    ( PHY_RXSYNC_HEADER ),   

         //  PHY Command
         .phy_txdetectrx_i       ( PHY_TXDETECTRX ),  
         .phy_txelecidle_i       ( PHY_TXELECIDLE ),                    
         .phy_txcompliance_i     ( PHY_TXCOMPLIANCE ), 
         .phy_rxpolarity_i       ( PHY_RXPOLARITY ),
         .phy_powerdown_i        ( PHY_POWERDOWN ), 
         .phy_rate_i             ( PHY_RATE ),

         .phy_txdetectrx_o       ( phy_txdetectrx_pl ),  
         .phy_txelecidle_o       ( phy_txelecidle_pl ),                    
         .phy_txcompliance_o     ( phy_txcompliance_pl ), 
         .phy_rxpolarity_o       ( phy_rxpolarity_pl ),
         .phy_powerdown_o        ( phy_powerdown_pl ), 
         .phy_rate_o             ( phy_rate_pl ),    

         //  PHY Status
         .phy_rxvalid_i          ( phy_rxvalid_pl ),
         .phy_phystatus_i        ( phy_phystatus_pl ),
         .phy_rxelecidle_i       ( phy_rxelecidle_pl ), 
         .phy_rxstatus_i         ( phy_rxstatus_pl ),

         .phy_rxvalid_o          ( PHY_RXVALID ),
         .phy_phystatus_o        ( PHY_PHYSTATUS ),
         .phy_rxelecidle_o       ( PHY_RXELECIDLE ), 
         .phy_rxstatus_o         ( PHY_RXSTATUS ),
        
         //  TX Driver
         .phy_txmargin_i         ( PHY_TXMARGIN ),          
         .phy_txswing_i          ( PHY_TXSWING ),           
         .phy_txdeemph_i         ( PHY_TXDEEMPH ),   

         .phy_txmargin_o         ( phy_txmargin_pl ),          
         .phy_txswing_o          ( phy_txswing_pl ),           
         .phy_txdeemph_o         ( phy_txdeemph_pl ),        

         //  TX Equalization (Gen3/4)
         .phy_txeq_ctrl_i        ( PHY_TXEQ_CTRL ),
         .phy_txeq_preset_i      ( PHY_TXEQ_PRESET ),
         .phy_txeq_coeff_i       ( PHY_TXEQ_COEFF ), 

         .phy_txeq_ctrl_o        ( phy_txeq_ctrl_pl ),
         .phy_txeq_preset_o      ( phy_txeq_preset_pl ),
         .phy_txeq_coeff_o       ( phy_txeq_coeff_pl ), 

         .phy_txeq_fs_i          ( phy_txeq_fs_pl ),           
         .phy_txeq_lf_i          ( phy_txeq_lf_pl ),           
         .phy_txeq_new_coeff_i   ( phy_txeq_new_coeff_pl ),
         .phy_txeq_done_i        ( phy_txeq_done_pl ),

         .phy_txeq_fs_o          ( PHY_TXEQ_FS ),           
         .phy_txeq_lf_o          ( PHY_TXEQ_LF ),           
         .phy_txeq_new_coeff_o   ( PHY_TXEQ_NEW_COEFF ),
         .phy_txeq_done_o        ( PHY_TXEQ_DONE ),   

         //  RX Equalization (Gen3/4)
         .phy_rxeq_ctrl_i        ( PHY_RXEQ_CTRL ), 
         .phy_rxeq_txpreset_i    ( PHY_RXEQ_TXPRESET ),

         .phy_rxeq_ctrl_o        ( phy_rxeq_ctrl_pl ), 
         .phy_rxeq_txpreset_o    ( phy_rxeq_txpreset_pl ),

         .phy_rxeq_preset_sel_i  ( phy_rxeq_preset_sel_pl ),
         .phy_rxeq_new_txcoeff_i ( phy_rxeq_new_txcoeff_pl ),
         .phy_rxeq_adapt_done_i  ( phy_rxeq_adapt_done_pl ),
         .phy_rxeq_done_i        ( phy_rxeq_done_pl ),

         .phy_rxeq_preset_sel_o  ( PHY_RXEQ_PRESET_SEL ),
         .phy_rxeq_new_txcoeff_o ( PHY_RXEQ_NEW_TXCOEFF ),
         .phy_rxeq_adapt_done_o  ( PHY_RXEQ_ADAPT_DONE ),
         .phy_rxeq_done_o        ( PHY_RXEQ_DONE ),

         // Assist Signals
         .as_mac_in_detect_i     ( AS_MAC_IN_DETECT ),
         .as_cdr_hold_req_i      ( AS_CDR_HOLD_REQ ),

         .as_mac_in_detect_o     ( as_mac_in_detect_pl ),
         .as_cdr_hold_req_o      ( as_cdr_hold_req_pl )
      );


         assign phy_txdetectrx_32b     = phy_txdetectrx_pl;
         assign phy_txelecidle_32b     = phy_txelecidle_pl;
         assign phy_txcompliance_32b   = phy_txcompliance_pl;
         assign phy_rxpolarity_32b     = phy_rxpolarity_pl;
         assign phy_powerdown_32b      = phy_powerdown_pl;
         assign phy_rate_32b           = phy_rate_pl;
         assign phy_txdata_64b         = phy_txdata_pl;
         assign phy_txdatak_32b        = phy_txdatak_pl;
         assign phy_txdata_valid_32b   = phy_txdata_valid_pl;
         assign phy_txstart_block_32b  = phy_txstart_block_pl;
         assign phy_txsync_header_32b  = phy_txsync_header_pl;
         assign phy_txeq_ctrl_pclk2    = phy_txeq_ctrl_pl;
         assign phy_txeq_preset_pclk2  = phy_txeq_preset_pl;
         assign phy_txeq_coeff_pclk2   = phy_txeq_coeff_pl;
         assign PHY_PCLK               = phy_pclk2;
         assign phy_rxdata_pl          = phy_rxdata_64b;          // 64b
         assign phy_rxdatak_pl         = phy_rxdatak_32b;
         assign phy_rxdata_valid_pl    = phy_rxdata_valid_32b;
         assign phy_rxstart_block_pl   = phy_rxstart_block_64b;   // 2b
         assign phy_rxsync_header_pl   = phy_rxsync_header_32b;
         assign phy_rxvalid_pl         = phy_rxvalid_pclk2;
         assign phy_phystatus_pl       = phy_phystatus_pclk2;
         assign PHY_PHYSTATUS_RST      = phy_phystatus_rst_pclk2;
         assign phy_rxstatus_raw       = phy_rxstatus_pclk2;
         assign phy_txeq_fs_pl         = phy_txeq_fs_pclk2;
         assign phy_txeq_lf_pl         = phy_txeq_lf_pclk2;
         assign phy_txeq_new_coeff_pl  = phy_txeq_new_coeff_pclk2;
         assign phy_txeq_done_pl       = phy_txeq_done_pclk2;
         assign phy_rxeq_preset_sel_pl = phy_rxeq_preset_sel_pclk2;
         assign phy_rxeq_new_txcoeff_pl= phy_rxeq_new_txcoeff_pclk2;
         assign phy_rxeq_done_pl       = phy_rxeq_done_pclk2;
         assign phy_rxeq_adapt_done_pl = phy_rxeq_adapt_done_pclk2;

 

   //--------------------------------------------------------------------------
   //  CDRHOLD Logic
   //--------------------------------------------------------------------------  

   `PHYREG(phy_pclk2, phy_phystatus_rst_pclk2, phy_rxelecidle_ff, phy_rxelecidle_pl[0], 'd1)
   `PHYREG(phy_pclk2, phy_phystatus_rst_pclk2, phy_rxelecidle_ff2, phy_rxelecidle_ff, 'd1)

   always @(*) begin 
      if (as_cdr_hold_req_pl & phy_rxelecidle_pl[0]) begin
         phy_rxcdrhold_wire   = 1'b1;
      end else if (phy_rxelecidle_ff2 & ~phy_rxelecidle_pl[0]) begin
         phy_rxcdrhold_wire   = 1'b0;
      end else begin
         phy_rxcdrhold_wire   = phy_rxcdrhold_pclk2;
      end
   end

   `PHYREG(phy_pclk2, phy_phystatus_rst_pclk2, phy_rxcdrhold_pclk2, phy_rxcdrhold_wire, 'd0)

   //--------------------------------------------------------------------------
   // Mask invalid RXSTATUS for Gen1/2 after EIOS, can be removed once GT fixes it
   //--------------------------------------------------------------------------

   assign phy_rxstatus_pl = phy_rxstatus_raw;


   //--------------------------------------------------------------------------
   //  UltraScale GTH PHY Wrapper
   //--------------------------------------------------------------------------   

   wire [((((PHY_LANE-1)>>2)+1)*16)-1:0]  gtcom_drpaddr_tie_off   = 'd0;
   wire [(PHY_LANE-1)>>2:0]               gtcom_drpen_tie_off     = 'd0;
   wire [(PHY_LANE-1)>>2:0]               gtcom_drpwe_tie_off     = 'd0;
   wire [((((PHY_LANE-1)>>2)+1)*16)-1:0]  gtcom_drpdi_tie_off     = 'd0;

   assign PHY_USERCLK   = ((PHY_USERCLK_FREQ == 3 && PHY_CORECLK_FREQ == 1) ||
                           (PHY_USERCLK_FREQ == 4 && PHY_CORECLK_FREQ == 2))  ? PHY_CORECLK : phy_userclk_int;

   assign PHY_MCAPCLK   = ((PHY_MCAPCLK_FREQ == 1 && PHY_USERCLK_FREQ == 1) ||
                           (PHY_MCAPCLK_FREQ == 2 && PHY_USERCLK_FREQ == 2))  ? phy_userclk_int : phy_mcapclk_int;

   generate
      if (FPGA_FAMILY == "USM") begin: diablo_gt
         xp4_usp_smsw_gt_phy_wrapper #(
            // Parameters
            .PHY_SIM_EN       ( PHY_SIM_EN ),     
            .PHY_GT_XCVR      ( (FPGA_XCVR == "Y")? "GTY": "GTH" ),
            .PHY_REFCLK_MODE  ( (PHY_ASYNC_EN == "FALSE")? 0: 1 ),
            .PHY_LANE         ( PHY_LANE ),   
            .PHY_MAX_SPEED    ( PHY_MAX_SPEED ),                    
            .PHY_REFCLK_FREQ  ( PHY_REFCLK_FREQ ),           
            .PHY_CORECLK_FREQ ( PHY_CORECLK_FREQ ),       
            .PHY_USERCLK_FREQ ( PHY_USERCLK_FREQ ),   
            .PHY_MCAPCLK_FREQ ( PHY_MCAPCLK_FREQ ),
            .PHY_GT_TXPRESET  ( PHY_GT_TXPRESET ),
            .PHY_LP_TXPRESET  ( PHY_LP_TXPRESET )
         ) diablo_gt_phy_wrapper_smsw (                                         
            // Clock & Reset Ports
            .PHY_REFCLK             ( PHY_REFCLK ),      
            .PHY_GTREFCLK           ( PHY_GTREFCLK ),               
            .PHY_RST_N              ( PHY_RST_N ),  
      
            .PHY_PCLK               ( phy_pclk2 ),  
            .PHY_PCLK2              ( phy_pclk ),  
            .PHY_CORECLK            ( PHY_CORECLK ), 
            .PHY_USERCLK            ( phy_userclk_int ),                          
            .PHY_MCAPCLK            ( phy_mcapclk_int ), // New in Diablo
                                                     
            // Serial Line Ports
            .PHY_RXP                ( PHY_RXP ),               
            .PHY_RXN                ( PHY_RXN ),               
                               
            .PHY_TXP                ( PHY_TXP ),               
            .PHY_TXN                ( PHY_TXN ),   
                                                                             
            // TX Data Ports 
            .PHY_TXDATA             ( phy_txdata_64b ),            
            .PHY_TXDATAK            ( phy_txdatak_32b ),                
            .PHY_TXDATA_VALID       ( phy_txdata_valid_32b ),                
            .PHY_TXSTART_BLOCK      ( phy_txstart_block_32b ),                      
            .PHY_TXSYNC_HEADER      ( phy_txsync_header_32b ),                                          
      
            // RX Data Ports 
            .PHY_RXDATA             ( phy_rxdata_64b ),            
            .PHY_RXDATAK            ( phy_rxdatak_32b ),                
            .PHY_RXDATA_VALID       ( phy_rxdata_valid_32b ),                
            .PHY_RXSTART_BLOCK      ( phy_rxstart_block_64b ),                      
            .PHY_RXSYNC_HEADER      ( phy_rxsync_header_32b ),                                          
      
            // PHY Command Port
            .PHY_TXDETECTRX         ( phy_txdetectrx_32b ),
            .PHY_TXELECIDLE         ( phy_txelecidle_32b ),                    
            .PHY_TXCOMPLIANCE       ( phy_txcompliance_32b ),                          
            .PHY_RXPOLARITY         ( phy_rxpolarity_32b ),            
            .PHY_POWERDOWN          ( phy_powerdown_32b ),
            .PHY_RATE               ( phy_rate_32b ),  
            .PHY_RXCDRHOLD          ( phy_rxcdrhold_pclk2 ),
          
            // PHY Status Ports
            .PHY_RXVALID            ( phy_rxvalid_pclk2 ),            
            .PHY_PHYSTATUS          ( phy_phystatus_pclk2 ),            
      
            .PHY_PHYSTATUS_RST      ( phy_phystatus_rst_pclk2 ),
            .PHY_RXELECIDLE         ( phy_rxelecidle_pl ),                    
            .PHY_RXSTATUS           ( phy_rxstatus_pclk2 ),                                            
          
            // TX Driver Ports
            .PHY_TXMARGIN           ( phy_txmargin_pl ),          
            .PHY_TXSWING            ( phy_txswing_pl ),   
            .PHY_TXDEEMPH           ( {1'b0, phy_txdeemph_pl} ),  // 2b in Diablo   
      
            // TX Equalization Ports for Gen3
            .PHY_TXEQ_CTRL          ( phy_txeq_ctrl_pclk2 ),
            .PHY_TXEQ_PRESET        ( phy_txeq_preset_pclk2 ),
            .PHY_TXEQ_COEFF         ( phy_txeq_coeff_pclk2 ),
      
            .PHY_TXEQ_FS            ( phy_txeq_fs_pclk2 ),           
            .PHY_TXEQ_LF            ( phy_txeq_lf_pclk2 ),           
            .PHY_TXEQ_NEW_COEFF     ( phy_txeq_new_coeff_pclk2 ),
            .PHY_TXEQ_DONE          ( phy_txeq_done_pclk2 ),
                                                                       
            // RX Equalization Ports for Gen3
            .PHY_RXEQ_CTRL          ( phy_rxeq_ctrl_pl ), 
            .PHY_RXEQ_PRESET        ( {PHY_LANE{3'b0}} ), 
            .PHY_RXEQ_LFFS          ( {PHY_LANE{6'b0}} ),         
            .PHY_RXEQ_TXPRESET      ( phy_rxeq_txpreset_pl ),
      
            .PHY_RXEQ_LFFS_SEL      ( phy_rxeq_preset_sel_pclk2 ),      
            .PHY_RXEQ_NEW_TXCOEFF   ( phy_rxeq_new_txcoeff_pclk2 ),   
            .PHY_RXEQ_DONE          ( phy_rxeq_done_pclk2 ),        
            .PHY_RXEQ_ADAPT_DONE    ( phy_rxeq_adapt_done_pclk2 ),
      
            // USB Ports
            .USB_TXONESZEROS        ( {PHY_LANE{1'b0}} ),   // New in Diablo
            .USB_RXEQTRAINING       ( {PHY_LANE{1'b0}} ),   // New in Diablo
            .USB_RXTERMINATION      ( {PHY_LANE{1'b0}} ),   // New in Diablo
            .USB_POWERPRESENT       ( ),  // New in Diablo
      
            // DRP Port
            .GT_DRPCLK              ( 1'b0 ),   // New in Diablo
            .GTCOM_DRPADDR          ( gtcom_drpaddr_tie_off ), // New in Diablo
            .GTCOM_DRPEN            ( gtcom_drpen_tie_off ),   // New in Diablo
            .GTCOM_DRPWE            ( gtcom_drpwe_tie_off ),   // New in Diablo
            .GTCOM_DRPDI            ( gtcom_drpdi_tie_off ),   // New in Diablo
            .GTCOM_DRPRDY           ( ),  // New in Diablo
            .GTCOM_DRPDO            ( ),  // New in Diablo 

            // Debug Ports   // Not used
            .DBG_RATE_DONE          ( {PHY_LANE{1'b0}} ),
            .DBG_RATE_START         ( ),  // New in Diablo
            .DBG_RATE_IDLE          ( ),  // New in Diablo
            .DBG_RXCDRLOCK          ( ),  // New in Diablo
            .DBG_GEN34_EIOS_DET     ( ),  // New in Diablo
            .DBG_TXOUTCLK           ( ),  // New in Diablo
            .DBG_RXOUTCLK           ( ),  // New in Diablo
            .DBG_TXOUTCLKFABRIC     ( ),  // New in Diablo
            .DBG_RXOUTCLKFABRIC     ( ),  // New in Diablo
            .DBG_TXOUTCLKPCS        ( ),  // New in Diablo
            .DBG_RXOUTCLKPCS        ( ),  // New in Diablo
            .DBG_RXRECCLKOUT        ( ),  // New in Diablo
            .DBG_TXPMARESET         ( {PHY_LANE{1'b0}} ),   // New in Diablo
            .DBG_RXPMARESET         ( {PHY_LANE{1'b0}} ),   // New in Diablo
            .DBG_TXPCSRESET         ( {PHY_LANE{1'b0}} ),   // New in Diablo
            .DBG_RXPCSRESET         ( {PHY_LANE{1'b0}} ),   // New in Diablo
            .DBG_RXBUFRESET         ( {PHY_LANE{1'b0}} ),   // New in Diablo
            .DBG_RXCDRRESET         ( {PHY_LANE{1'b0}} ),   // New in Diablo
            .DBG_RXDFELPMRESET      ( {PHY_LANE{1'b0}} ),   // New in Diablo
            .DBG_RRST_N             ( ),  // New in Diablo
            .DBG_PRST_N             ( ),  // New in Diablo
            .DBG_GTPOWERGOOD        ( ),  // New in Diablo
            .DBG_CPLLLOCK           ( ),  // New in Diablo
            .DBG_QPLL0LOCK          ( ),  // New in Diablo
            .DBG_QPLL1LOCK          ( ),  // New in Diablo
            .DBG_TXPROGDIVRESETDONE ( ),  // New in Diablo
            .DBG_TXPMARESETDONE     ( ),  // New in Diablo
            .DBG_RXPMARESETDONE     ( ),  // New in Diablo
            .DBG_TXRESETDONE        ( ),  // New in Diablo
            .DBG_RXRESETDONE        ( ),  // New in Diablo
            .DBG_TXSYNCDONE         ( ),  // New in Diablo
            .DBG_RST_IDLE           ( ),  // New in Diablo
      
            // PRBS Debug Ports
            .DBG_LOOPBACK           ( 3'b0 ),   // New in Diablo
            .DBG_PRBSSEL            ( 4'b0 ),   // New in Diablo
            .DBG_TXPRBSFORCEERR     ( 1'b0 ),   // New in Diablo
            .DBG_RXPRBSCNTRESET     ( 1'b0 ),   // New in Diablo
            .DBG_RXPRBSERR          ( ),  // New in Diablo
            .DBG_RXPRBSLOCKED       ( ),  // New in Diablo
            .PHY_PCIE_MAC_IN_DETECT ( as_mac_in_detect_pl ) // New in Diablo
         );
      end 
   endgenerate

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_gt_phy_wrapper.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
//  Design  :  Diablo PHY Wrapper REFERENCE DESIGN
//  Module  :  PHY Wrapper Top
//--------------------------------------------------------------------------------------------------
//  *** XILINX INTERNAL *** 
//--------------------------------------------------------------------------------------------------
//  Version :  0.73
//--------------------------------------------------------------------------------------------------

//--------------------------------------------------------------------------------------------------
//  PHY Wrapper Design Hierarchy in Static Mode
//--------------------------------------------------------------------------------------------------
//  PHY Wrapper Top :
//      - Clock 
//      - Reset
//      - PHY Lane :
//          - TX Equalization (Gen3/Gen4)
//          - RX Equalization (Gen3/Gen4)
//          - GT Channel (one channel for every lane)
//      - PHY Quad :
//          - GT Common (one quad for every four lanes)
//--------------------------------------------------------------------------------------------------

//--------------------------------------------------------------------------------------------------
//  PHY Wrapper Design Hierarchy in GT Wizard Mode
//--------------------------------------------------------------------------------------------------
//  PHY Wrapper Top :
//      - Clock 
//      - Reset
//      - PHY Lane :
//          - TX Equalization (Gen3/Gen4)
//          - RX Equalization (Gen3/Gen4)
//      - GT Wizard Top :
//          - GT Wizard Core
//              - GT Channel (one channel for every lane)
//              - GT Common (one quad for every four lanes)
//--------------------------------------------------------------------------------------------------

//--------------------------------------------------------------------------------------------------
//  PHY Wrapper User Parameter Encoding
//--------------------------------------------------------------------------------------------------
//  PHY_SIM_EN                : "FALSE" = Normal
//                            : "TRUE"  = Simulation
//  PHY_GT_XCVR               : "GTH" = GTH Transceiver
//                            : "GTY" = GTY Transceiver
//                            : "GTY64" = GTY with 64-bit support for PCIe Gen4
//  PHY_MODE                  : 0 = PCIe 4.0
//                            : 1 = USB  3.0
//  PHY_REFCLK_MODE           : 0 =          0 ppm (Common   REFCLK)
//                            : 1 = up to  600 ppm (Seperate REFCLK without SSC)
//                            : 2 = up to 5600 ppm (Seperate REFCLK with independent SSC)
//  PHY_GTWIZARD              : "FALSE" = Use Static Wrapper mode
//                            : "TRUE"  = Use GT Wizard Generated Wrapper mode
//  PHY_LANE                  : 1, 2, 4, 8, 16 
//  PHY_MAX_SPEED             : 1 = PCIe Gen1 ( 2.5 Gbps) Capable or USB3 Gen1 ( 5.0 Gb/s)        
//                            : 2 = PCIe Gen2 ( 5.0 Gbps) Capable
//                            : 3 = PCIe Gen3 ( 8.0 Gbps) Capable 
//                            : 4 = PCIe Gen4 (16.0 Gbps) Capable
//  PHY_GEN12_CDR_CTRL_ON_EIDLE : "FALSE" = Will not auto reset CDR upon EIOS detection (Gen1/Gen2)
//                            : "TRUE"  = Will     auto reset CDR upon EIOS detection (Gen1/Gen2)
//  PHY_GEN34_CDR_CTRL_ON_EIDLE : "FALSE" = Will not auto reset CDR upon EIOS detection (Gen3/Gen4)
//                            : "TRUE"  = Will     auto reset CDR upon EIOS detection (Gen3/Gen4)
//  PHY_REFCLK_FREQ           : 0 = 100.0 MHz 
//                            : 1 = 125.0 MHz
//                            : 2 = 250.0 MHz
//  PHY_CORECLK_FREQ          : 1 = 250.0 MHz
//                            : 2 = 500.0 MHz
//  PHY_USERCLK_FREQ          : 1 =  62.5 MHz
//                            : 2 = 125.0 MHz
//                            : 3 = 250.0 MHz
//                            : 4 = 500.0 MHz
//  PHY_MCAPCLK_FREQ          : 1 =  62.5 MHz
//                            : 2 = 125.0 MHz
//                            : 3 = 250.0 MHz
//                            : 4 = 500.0 MHz
//  PHY_GT_TXPRESET           : 0 to 10 
//  PHY_LP_TXPRESET           : 0 to 10 
//--------------------------------------------------------------------------------------------------

`timescale 1ps / 1ps

//--------------------------------------------------------------------------------------------------
//  PHY Wrapper Top
//--------------------------------------------------------------------------------------------------
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_gt_phy_wrapper #
(
    //--------------------------------------------------------------------------
    //  Parameters
    //--------------------------------------------------------------------------
    parameter         PHY_SIM_EN                 = "FALSE",   
    parameter         PHY_GT_XCVR                = "GTY",
    parameter         PHY_GTWIZARD               = "FALSE",
    parameter integer PHY_MODE                   = 0,  
    parameter integer PHY_REFCLK_MODE            = 0,       
    parameter integer PHY_LANE                   = 1,   
    parameter integer PHY_MAX_SPEED              = 4,  
    parameter         PHY_GEN12_CDR_CTRL_ON_EIDLE = "TRUE",                
    parameter         PHY_GEN34_CDR_CTRL_ON_EIDLE = "TRUE",     
    parameter integer PHY_REFCLK_FREQ            = 0, 
    parameter integer PHY_CORECLK_FREQ           = 2,       
    parameter integer PHY_USERCLK_FREQ           = 4,           
    parameter integer PHY_MCAPCLK_FREQ           = 4,    
    parameter integer PHY_GT_TXPRESET            = 0,
    parameter integer PHY_LP_TXPRESET            = 4         
)                                                            
(                                         
    //--------------------------------------------------------------------------
    //  Clock & Reset Ports
    //--------------------------------------------------------------------------
    input                               PHY_REFCLK,                             // For PHY Wrapper
    input                               PHY_GTREFCLK,                           // For GT
    input                               PHY_RST_N,                              // System RST
   
    output                              PHY_PCLK,                               
    output                              PHY_PCLK2,                              // For PCIe IP                          
    output                              PHY_CORECLK,                            // For PCIe IP
    output                              PHY_USERCLK,                            // For PCIe IP
    output                              PHY_MCAPCLK,                            // For PCIe IP
  
    //--------------------------------------------------------------------------
    //  Serial Line Ports
    //--------------------------------------------------------------------------
    input       [PHY_LANE-1:0]          PHY_RXP,               
    input       [PHY_LANE-1:0]          PHY_RXN,               

    output      [PHY_LANE-1:0]          PHY_TXP,               
    output      [PHY_LANE-1:0]          PHY_TXN,   
 
    //--------------------------------------------------------------------------
    //  TX Data Ports 
    //--------------------------------------------------------------------------
    input       [(PHY_LANE*64)-1:0]     PHY_TXDATA,         
    input       [(PHY_LANE* 2)-1:0]     PHY_TXDATAK,    
    input       [PHY_LANE-1:0]          PHY_TXDATA_VALID,
    input       [PHY_LANE-1:0]          PHY_TXSTART_BLOCK,      
    input       [(PHY_LANE* 2)-1:0]     PHY_TXSYNC_HEADER,                    

    //--------------------------------------------------------------------------
    //  RX Data Ports 
    //--------------------------------------------------------------------------
    output      [(PHY_LANE*64)-1:0]     PHY_RXDATA,         
    output      [(PHY_LANE* 2)-1:0]     PHY_RXDATAK,       
    output      [PHY_LANE-1:0]          PHY_RXDATA_VALID,         
    output      [(PHY_LANE* 2)-1:0]     PHY_RXSTART_BLOCK,  
    output      [(PHY_LANE* 2)-1:0]     PHY_RXSYNC_HEADER,
    
    //--------------------------------------------------------------------------
    //  PHY Command Port
    //--------------------------------------------------------------------------
    input                               PHY_TXDETECTRX,        
    input       [PHY_LANE-1:0]          PHY_TXELECIDLE,        
    input       [PHY_LANE-1:0]          PHY_TXCOMPLIANCE,      
    input       [PHY_LANE-1:0]          PHY_RXPOLARITY,        
    input       [1:0]                   PHY_POWERDOWN,         
    input       [1:0]                   PHY_RATE,    
    input                               PHY_RXCDRHOLD,                          // For Gen3/Gen4 RX EQ             
    
    //--------------------------------------------------------------------------   
    //  PHY Status Ports
    //-------------------------------------------------------------------------- 
    output      [PHY_LANE-1:0]          PHY_RXVALID,               
    output      [PHY_LANE-1:0]          PHY_PHYSTATUS,          
    output                              PHY_PHYSTATUS_RST,                      // For PCIe IP
    output      [PHY_LANE-1:0]          PHY_RXELECIDLE,         
    output      [(PHY_LANE*3)-1:0]      PHY_RXSTATUS,                       
    
    //--------------------------------------------------------------------------
    //  TX Driver Ports
    //--------------------------------------------------------------------------
    input       [ 2:0]                  PHY_TXMARGIN,          
    input                               PHY_TXSWING,           
    input       [ 1:0]                  PHY_TXDEEMPH,    
    
    //--------------------------------------------------------------------------   
    //  TX Equalization Ports (Gen3/Gen4)
    //--------------------------------------------------------------------------  
    input       [(PHY_LANE*2)-1:0]      PHY_TXEQ_CTRL,      
    input       [(PHY_LANE*4)-1:0]      PHY_TXEQ_PRESET,       
    input       [(PHY_LANE*6)-1:0]      PHY_TXEQ_COEFF,                                                            

    output      [ 5:0]                  PHY_TXEQ_FS,           
    output      [ 5:0]                  PHY_TXEQ_LF,           
    output      [(PHY_LANE*18)-1:0]     PHY_TXEQ_NEW_COEFF,        
    output      [PHY_LANE-1:0]          PHY_TXEQ_DONE,         

    //--------------------------------------------------------------------------
    //  RX Equalization Ports (Gen3/Gen4)
    //--------------------------------------------------------------------------                                                
    input       [(PHY_LANE*2)-1:0]      PHY_RXEQ_CTRL,     
    input       [(PHY_LANE*3)-1:0]      PHY_RXEQ_PRESET,  
    input       [(PHY_LANE*4)-1:0]      PHY_RXEQ_TXPRESET,      
    input       [(PHY_LANE*6)-1:0]      PHY_RXEQ_LFFS,                                                         

    output      [PHY_LANE-1:0]          PHY_RXEQ_LFFS_SEL,    
    output      [(PHY_LANE*18)-1:0]     PHY_RXEQ_NEW_TXCOEFF,   
    output      [PHY_LANE-1:0]          PHY_RXEQ_ADAPT_DONE,     
    output      [PHY_LANE-1:0]          PHY_RXEQ_DONE,         
    
    //--------------------------------------------------------------------------
    //  GT Channel Ports (USB3)
    //--------------------------------------------------------------------------
    input       [PHY_LANE-1:0]          USB_TXONESZEROS,                        
    input       [PHY_LANE-1:0]          USB_RXEQTRAINING,                       
    input       [PHY_LANE-1:0]          USB_RXTERMINATION,                        
    
    output      [PHY_LANE-1:0]          USB_POWERPRESENT,    
    
    //--------------------------------------------------------------------------
    //  GT Common DRP Ports 
    //--------------------------------------------------------------------------
    input                                           GT_DRPCLK,
    input       [((((PHY_LANE-1)>>2)+1)*16)-1:0]    GTCOM_DRPADDR,                                       
    input       [   (PHY_LANE-1)>>2          :0]    GTCOM_DRPEN,                                             
    input       [   (PHY_LANE-1)>>2          :0]    GTCOM_DRPWE,     
    input       [((((PHY_LANE-1)>>2)+1)*16)-1:0]    GTCOM_DRPDI,                                      
                                                                         
    output      [   (PHY_LANE-1)>>2          :0]    GTCOM_DRPRDY,    
    output      [((((PHY_LANE-1)>>2)+1)*16)-1:0]    GTCOM_DRPDO,       
    
    //----------------------------------------------------------------------------------------------
    //  GT Debug Ports
    //----------------------------------------------------------------------------------------------       
    input       [PHY_LANE-1:0]          DBG_RATE_DONE,
    
    output      [PHY_LANE-1:0]          DBG_RATE_START,             
    output      [PHY_LANE-1:0]          DBG_RATE_IDLE,
    output      [PHY_LANE-1:0]          DBG_RXCDRLOCK,     
    output      [PHY_LANE-1:0]          DBG_GEN34_EIOS_DET, 
    
    //--------------------------------------------------------------------------
    // CLK Debug Ports (Requires BUFG if used)
    //--------------------------------------------------------------------------
    output      [PHY_LANE-1:0]          DBG_TXOUTCLK, 
    output      [PHY_LANE-1:0]          DBG_RXOUTCLK, 
    output      [PHY_LANE-1:0]          DBG_TXOUTCLKFABRIC,                                                              
    output      [PHY_LANE-1:0]          DBG_RXOUTCLKFABRIC,                                                              
    output      [PHY_LANE-1:0]          DBG_TXOUTCLKPCS,                                                              
    output      [PHY_LANE-1:0]          DBG_RXOUTCLKPCS,                 
    output      [PHY_LANE-1:0]          DBG_RXRECCLKOUT, 
        
    //--------------------------------------------------------------------------
    // RST Debug Ports
    //--------------------------------------------------------------------------     
    input       [PHY_LANE-1:0]          DBG_TXPMARESET,                                            
    input       [PHY_LANE-1:0]          DBG_RXPMARESET,                                            
    input       [PHY_LANE-1:0]          DBG_TXPCSRESET,   
    input       [PHY_LANE-1:0]          DBG_RXPCSRESET,
    input       [PHY_LANE-1:0]          DBG_RXBUFRESET,
    input       [PHY_LANE-1:0]          DBG_RXCDRRESET,
    input       [PHY_LANE-1:0]          DBG_RXDFELPMRESET,
   
    output                              DBG_RRST_N,
    output                              DBG_PRST_N,       
    output      [PHY_LANE-1:0]          DBG_GTPOWERGOOD,  
    output      [PHY_LANE-1:0]          DBG_CPLLLOCK,      
    output      [(PHY_LANE-1)>>2:0]     DBG_QPLL0LOCK,    
    output      [(PHY_LANE-1)>>2:0]     DBG_QPLL1LOCK,  
    output      [PHY_LANE-1:0]          DBG_TXPROGDIVRESETDONE,
    output      [PHY_LANE-1:0]          DBG_TXPMARESETDONE,   
    output      [PHY_LANE-1:0]          DBG_RXPMARESETDONE, 
    output      [PHY_LANE-1:0]          DBG_TXRESETDONE,
    output      [PHY_LANE-1:0]          DBG_RXRESETDONE,    
    output      [PHY_LANE-1:0]          DBG_TXSYNCDONE,  
    output                              DBG_RST_IDLE,               

    //--------------------------------------------------------------------------
    //  PRBS Debug Ports
    //--------------------------------------------------------------------------
    input       [ 2:0]                  DBG_LOOPBACK,                                              
    input       [ 3:0]                  DBG_PRBSSEL,
    input                               DBG_TXPRBSFORCEERR,
    input                               DBG_RXPRBSCNTRESET,                                                                                                      

    output      [PHY_LANE-1:0]          DBG_RXPRBSERR,                                              
    output      [PHY_LANE-1:0]          DBG_RXPRBSLOCKED,
    
    //---------------------------------------------------------------------------
    //   Receiver Detect (Remote TX detecting our RX)
    //---------------------------------------------------------------------------
    input                               PHY_PCIE_MAC_IN_DETECT 
);

//--------------------------------------------------------------------------------------------------
//  Internal Signals
//--------------------------------------------------------------------------------------------------

    //--------------------------------------------------------------------------
    //  Clock 
    //--------------------------------------------------------------------------
    wire                                pclk; 
    wire                                pclk2_gt;
  
    //--------------------------------------------------------------------------
    //  Reset
    //--------------------------------------------------------------------------
    wire                                rrst_n;
    wire                                prst_n;
    
    wire                                rst_cpllpd;
    wire                                rst_cpllreset;  
    wire                                rst_qpllpd;  
    wire                                rst_qpllreset;
    wire                                rst_txprogdivreset;
    wire                                rst_gtreset;
    wire                                rst_userrdy; 
    wire                                rst_txsync_start;
    wire                                rst_idle;

    //--------------------------------------------------------------------------
    //  TX Equalization (Gen3/Gen4)
    //-------------------------------------------------------------------------- 
    wire        [(PHY_LANE*5)-1:0]      txeq_precursor; 
    wire        [(PHY_LANE*7)-1:0]      txeq_maincursor; 
    wire        [(PHY_LANE*5)-1:0]      txeq_postcursor; 
    wire        [(PHY_LANE*18)-1:0]     txeq_new_coeff; 
    wire        [PHY_LANE-1:0]          txeq_done;  
    
    //--------------------------------------------------------------------------
    //  RX Equalization (Gen3/Gen4)
    //-------------------------------------------------------------------------- 
    wire        [PHY_LANE-1:0]          rxeq_lffs_sel;   
    wire        [(PHY_LANE*18)-1:0]     rxeq_new_txcoeff;    
    wire        [PHY_LANE-1:0]          rxeq_adapt_done;     
    wire        [PHY_LANE-1:0]          rxeq_done;   
    
    //--------------------------------------------------------------------------
    //  GT Channel 
    //--------------------------------------------------------------------------
    wire        [PHY_LANE-1:0]          gt_bufgtce;    
    wire        [(PHY_LANE*3)-1:0]      gt_bufgtcemask;
    wire        [PHY_LANE-1:0]          gt_bufgtreset;
    wire        [(PHY_LANE*3)-1:0]      gt_bufgtrstmask;   
    wire        [(PHY_LANE*9)-1:0]      gt_bufgtdiv;
    wire        [PHY_LANE-1:0]          gt_txoutclk; 

    wire        [PHY_LANE-1:0]          gt_gtpowergood;
    wire        [PHY_LANE-1:0]          gt_txprogdivresetdone;
    wire        [PHY_LANE-1:0]          gt_txresetdone;
    wire        [PHY_LANE-1:0]          gt_rxresetdone;
    
    wire        [(PHY_LANE*3)-1:0]      gt_qpllrate;                           
    
    wire        [PHY_LANE-1:0]          gt_phystatus;
    wire        [PHY_LANE-1:0]          gt_rxelecidle;
    
    wire        [PHY_LANE-1:0]          gt_pcieuserphystatusrst;
    wire        [(PHY_LANE*2)-1:0]      gt_pcierateqpllpd;                 
    wire        [(PHY_LANE*2)-1:0]      gt_pcierateqpllreset;               
    wire        [PHY_LANE-1:0]          gt_pcierateidle;            
    wire        [PHY_LANE-1:0]          gt_pciesynctxsyncdone;                 
    wire        [PHY_LANE-1:0]          gt_pcierategen3;  
    wire        [PHY_LANE-1:0]          gt_pcieusergen3rdy; 
    wire        [PHY_LANE-1:0]          gt_pcieuserratestart;  
    
    wire        [PHY_LANE-1:0]          gt_txphaligndone;                                          
    wire        [PHY_LANE-1:0]          gt_txsyncout;                          
    
    wire        [PHY_LANE-1:0]          gt_cplllock;     
    wire        [PHY_LANE-1:0]          gt_rxcdrlock;    
    
    wire        [PHY_LANE-1:0]          gt_rxcdrhold;
    wire        [PHY_LANE-1:0]          gt_gen34_eios_det;
                                   
    wire        [PHY_LANE-1:0]          gt_rxratedone;
    wire        [PHY_LANE-1:0]          gt_rxtermination;

    //--------------------------------------------------------------------------
    //  GT Common
    //--------------------------------------------------------------------------
    wire        [(PHY_LANE-1)>>2:0]     gtcom_qpll0lock;
    wire        [(PHY_LANE-1)>>2:0]     gtcom_qpll0outclk;          
    wire        [(PHY_LANE-1)>>2:0]     gtcom_qpll0outrefclk;       
                                       
    wire        [(PHY_LANE-1)>>2:0]     gtcom_qpll1lock;
    wire        [(PHY_LANE-1)>>2:0]     gtcom_qpll1outclk;          
    wire        [(PHY_LANE-1)>>2:0]     gtcom_qpll1outrefclk;       

    //--------------------------------------------------------------------------
    //  Signals for GT Common
    //--------------------------------------------------------------------------
    wire        [(PHY_LANE-1)>>2:0]     qpll0pd;                    
    wire        [(PHY_LANE-1)>>2:0]     qpll0reset;                 
    wire        [(PHY_LANE-1)>>2:0]     qpll1pd;                    
    wire        [(PHY_LANE-1)>>2:0]     qpll1reset;                 
                                       
    //--------------------------------------------------------------------------
    //  Signals converted from per lane
    //--------------------------------------------------------------------------
    wire                                qpll0lock_all;                         
    wire                                qpll1lock_all;
    wire                                txsyncallin_all;                       

    //--------------------------------------------------------------------------
    //  GT DRP signals
    //--------------------------------------------------------------------------    
    
    wire        [(PHY_LANE*10)-1:0]     gt_drpaddr = {PHY_LANE{10'd0}}; 
    wire        [PHY_LANE-1:0]          gt_drpen   = {PHY_LANE{1'b0}};
    wire        [PHY_LANE-1:0]          gt_drpwe   = {PHY_LANE{1'b0}};
    wire        [(PHY_LANE*16)-1:0]     gt_drpdi   = {PHY_LANE{16'd0}};

    wire        [PHY_LANE-1:0]          gt_drprdy;
    wire        [(PHY_LANE*16)-1:0]     gt_drpdo;  

    //--------------------------------------------------------------------------
    // Reciever Detect RX termination signals 
    //--------------------------------------------------------------------------    
    
    wire        [PHY_LANE-1:0]         rxterm_rxtermination;

    //--------------------------------------------------------------------------
    //  CDR Control signals
    //-------------------------------------------------------------------------- 
    
    wire        [PHY_LANE-1:0]         cdrctrl_rxcdrhold;
    wire        [PHY_LANE-1:0]         cdrctrl_rxcdrfreqreset;
    wire        [PHY_LANE-1:0]         cdrctrl_resetovrd;
    
    //--------------------------------------------------------------------------
    //  PHYSTATUS Reset Synchronizer for PCLK
    //--------------------------------------------------------------------------

    (* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO", keep = "true", max_fanout = 500 *) reg [3:0] rst_psrst_n_r;

    //----
    //  
    //----

    wire                                bufg_gt_ce;
    wire                                bufg_gt_reset;
   (* keep = "true" *) wire [2:0]       PHY_TXOUTCLKSEL;

    assign bufg_gt_ce = rrst_n ? gt_bufgtce[0] : 1'b1;
    assign bufg_gt_reset = !rst_cpllreset ? gt_bufgtreset[0] : 1'b0;
    assign PHY_TXOUTCLKSEL = rst_cpllreset ? 3'h3 : 3'h5; 

   // 64-bit support for PCIe Gen4
    localparam PHY_GEN4_64BIT_EN = (PHY_GT_XCVR == "GTY64") ? "TRUE" : "FALSE";
//--------------------------------------------------------------------------------------------------
//  PHY Clock 
//--------------------------------------------------------------------------------------------------
xp4_usp_smsw_gt_phy_clk #
(
    .PHY_MAX_SPEED                      (PHY_MAX_SPEED),
    .PHY_GEN4_64BIT_EN                  (PHY_GEN4_64BIT_EN),
    .PHY_CORECLK_FREQ                   (PHY_CORECLK_FREQ),   
    .PHY_USERCLK_FREQ                   (PHY_USERCLK_FREQ),  
    .PHY_MCAPCLK_FREQ                   (PHY_MCAPCLK_FREQ) 
)
phy_clk_smsw_i
(
    //--------------------------------------------------------------------------
    //  CLK Port
    //--------------------------------------------------------------------------
    .CLK_TXOUTCLK                       (gt_txoutclk[0]),                       // From master lane 0
    .CLK_PCLK2_GT                       (pclk2_gt),                             // To all [TX/RX]USRCLK2

    //--------------------------------------------------------------------------
    //  PCLK Ports
    //--------------------------------------------------------------------------   
    .CLK_PCLK_CE                        (bufg_gt_ce),                  
    .CLK_PCLK_CEMASK                    (gt_bufgtcemask[0]), 
    .CLK_PCLK_CLR                       (bufg_gt_reset),                     
    .CLK_PCLK_CLRMASK                   (gt_bufgtrstmask[0]),   
    .CLK_PCLK_DIV                       (gt_bufgtdiv[2:0]),    
    .CLK_PCLK                           (pclk),
    
    //--------------------------------------------------------------------------
    //  PCLK2 Ports
    //--------------------------------------------------------------------------    
    .CLK_PCLK2_CE                       (bufg_gt_ce),                  
    .CLK_PCLK2_CEMASK                   (gt_bufgtcemask[0]), 
    .CLK_PCLK2_CLR                      (bufg_gt_reset),                     
    .CLK_PCLK2_CLRMASK                  (gt_bufgtrstmask[0]),   
    .CLK_PCLK2_DIV                      (gt_bufgtdiv[8:6]),    
    .CLK_PCLK2                          (PHY_PCLK2),
    
    //--------------------------------------------------------------------------
    //  CORECLK Ports
    //--------------------------------------------------------------------------
    .CLK_CORECLK_CE                     (bufg_gt_ce),                               
    .CLK_CORECLK_CEMASK                 (rst_idle),            
    .CLK_CORECLK_CLR                    (bufg_gt_reset),                     
    .CLK_CORECLK_CLRMASK                (rst_idle),                                        
    .CLK_CORECLK                        (PHY_CORECLK), 
    
    //--------------------------------------------------------------------------
    //  USERCLK Ports
    //--------------------------------------------------------------------------                      
    .CLK_USERCLK_CE                     (bufg_gt_ce),                       
    .CLK_USERCLK_CEMASK                 (rst_idle),
    .CLK_USERCLK_CLR                    (bufg_gt_reset),                     
    .CLK_USERCLK_CLRMASK                (rst_idle),
    .CLK_USERCLK                        (PHY_USERCLK),
    
    //--------------------------------------------------------------------------
    //  MCAPCLK Ports
    //--------------------------------------------------------------------------                     
    .CLK_MCAPCLK_CE                     (bufg_gt_ce),
    .CLK_MCAPCLK_CEMASK                 (rst_idle),
    .CLK_MCAPCLK_CLR                    (bufg_gt_reset),                     
    .CLK_MCAPCLK_CLRMASK                (rst_idle),
    .CLK_MCAPCLK                        (PHY_MCAPCLK) 
);



//--------------------------------------------------------------------------------------------------
//  PHY Reset
//--------------------------------------------------------------------------------------------------
xp4_usp_smsw_gt_phy_rst #
(
    .PHY_LANE                           (PHY_LANE),
    .PHY_MAX_SPEED                      (PHY_MAX_SPEED)            
)
phy_rst_smsw_i
(
    //-------------------------------------------------------------------------- 
    //  Input Ports
    //--------------------------------------------------------------------------       
    .RST_REFCLK                         (PHY_REFCLK),   
    .RST_PCLK                           (pclk),                         
    .RST_N                              (PHY_RST_N),  
    .RST_GTPOWERGOOD                    (gt_gtpowergood),                
    .RST_CPLLLOCK                       (gt_cplllock),   
    .RST_QPLL1LOCK                      (gtcom_qpll1lock), 
    .RST_QPLL0LOCK                      (gtcom_qpll0lock),
    .RST_TXPROGDIVRESETDONE             (gt_txprogdivresetdone),                           
    .RST_TXRESETDONE                    (gt_txresetdone), 
    .RST_RXRESETDONE                    (gt_rxresetdone), 
    .RST_TXSYNC_DONE                    (gt_pciesynctxsyncdone),     
    .RST_PHYSTATUS                      (gt_phystatus),                                             

    //-------------------------------------------------------------------------- 
    //  Output Ports
    //--------------------------------------------------------------------------   
    .RST_RRST_N                         (rrst_n),
    .RST_PRST_N                         (prst_n), 
    .RST_CPLLPD                         (rst_cpllpd),               
    .RST_CPLLRESET                      (rst_cpllreset),  
    .RST_QPLLPD                         (rst_qpllpd),
    .RST_QPLLRESET                      (rst_qpllreset),  
    .RST_TXPROGDIVRESET                 (rst_txprogdivreset),                              
    .RST_GTRESET                        (rst_gtreset),               
    .RST_USERRDY                        (rst_userrdy),   
    .RST_TXSYNC_START                   (rst_txsync_start),                                
    .RST_IDLE                           (rst_idle)                          
);
   


//--------------------------------------------------------------------------------------------------
//  Generate PHY Lane - Begin
//--------------------------------------------------------------------------------------------------
genvar i;   
    
generate for (i=0; i<PHY_LANE; i=i+1) 

    begin : phy_lane
    
    //----------------------------------------------------------------------------------------------
    //  PHY TX Equalization (Gen3)
    //----------------------------------------------------------------------------------------------
    xp4_usp_smsw_gt_phy_txeq #
    (
        .PHY_GT_TXPRESET                (PHY_GT_TXPRESET)                
    )
    phy_txeq_smsw_i
    (
        //---------------------------------------------------------------------- 
        //  Input Ports
        //----------------------------------------------------------------------  
        .TXEQ_CLK                       (pclk),
        .TXEQ_RST_N                     (prst_n),    
        .TXEQ_CTRL                      (PHY_TXEQ_CTRL[(2*i)+1:(2*i)]), 
        .TXEQ_PRESET                    (PHY_TXEQ_PRESET[(4*i)+3:(4*i)]), 
        .TXEQ_COEFF                     (PHY_TXEQ_COEFF[(6*i)+5:(6*i)]),

        //---------------------------------------------------------------------- 
        //  Output Ports
        //----------------------------------------------------------------------   
        .TXEQ_PRECURSOR                 (txeq_precursor[(5*i)+4:(5*i)]),        
        .TXEQ_MAINCURSOR                (txeq_maincursor[(7*i)+6:(7*i)]),       
        .TXEQ_POSTCURSOR                (txeq_postcursor[(5*i)+4:(5*i)]),       
        .TXEQ_NEW_COEFF                 (txeq_new_coeff[(18*i)+17:(18*i)]),          
        .TXEQ_DONE                      (txeq_done[i])      
    );                                                   



    //----------------------------------------------------------------------------------------------
    //  PHY RX Equalization (Gen3)
    //----------------------------------------------------------------------------------------------
    xp4_usp_smsw_gt_phy_rxeq #
    (
        .PHY_SIM_EN                     (PHY_SIM_EN),
        .PHY_LP_TXPRESET                (PHY_LP_TXPRESET)                
    )
    phy_rxeq_smsw_i
    (
        //---------------------------------------------------------------------- 
        //  Input Ports
        //----------------------------------------------------------------------  
        .RXEQ_CLK                       (pclk),
        .RXEQ_RST_N                     (prst_n),  
        .RXEQ_CTRL                      (PHY_RXEQ_CTRL[(2*i)+1:(2*i)]), 
        .RXEQ_PRESET                    (PHY_RXEQ_PRESET[(3*i)+2:(3*i)]), 
        .RXEQ_TXPRESET                  (PHY_RXEQ_TXPRESET[(4*i)+3:(4*i)]),
        .RXEQ_TXCOEFF                   (PHY_TXEQ_COEFF[(6*i)+5:(6*i)]),
        .RXEQ_LFFS                      (PHY_RXEQ_LFFS[(6*i)+5:(6*i)]),

        //---------------------------------------------------------------------- 
        //  Output Ports
        //----------------------------------------------------------------------     
        .RXEQ_LFFS_SEL                  (rxeq_lffs_sel[i]),   
        .RXEQ_NEW_TXCOEFF               (rxeq_new_txcoeff[(18*i)+17:(18*i)]),    
        .RXEQ_ADAPT_DONE                (rxeq_adapt_done[i]),      
        .RXEQ_DONE                      (rxeq_done[i])      
    );

    //----------------------------------------------------------------------------------------------
    //  Receiver detect RX termination
    //----------------------------------------------------------------------------------------------    
    xp4_usp_smsw_gt_receiver_detect_rxterm #
    ( 
      .CONSECUTIVE_CYCLE_OF_RXELECIDLE ((PHY_REFCLK_FREQ==0)?64:(PHY_REFCLK_FREQ==1)?80:160)
    )
    receiver_detect_termination_smsw_i
    (
      //---------- Input -------------------------------------
      .RXTERM_CLK                        (PHY_REFCLK), 
      .RXTERM_RST_N                      (rrst_n), 
      .RXTERM_RXELECIDLE                 (PHY_RXELECIDLE[i]), 
      .RXTERM_MAC_IN_DETECT              (PHY_PCIE_MAC_IN_DETECT), 
    
      //---------- Output ------------------------------------
      .RXTERM_RXTERMINATION              (rxterm_rxtermination[i]),
      .RXTERM_FSM                        () 
    );
    
    assign gt_rxtermination[i] = (PHY_MODE == 0) ? rxterm_rxtermination[i] : USB_RXTERMINATION[i];

    //--------------------------------------------------------------------------------------------------
    //  Reset CDR upon EIOS/EIDLE detection
    //--------------------------------------------------------------------------------------------------
    xp4_usp_smsw_gt_cdr_ctrl_on_eidle #
    (
        .PHY_GEN12_CDR_CTRL_ON_EIDLE (PHY_GEN12_CDR_CTRL_ON_EIDLE),   
        .PHY_GEN34_CDR_CTRL_ON_EIDLE (PHY_GEN34_CDR_CTRL_ON_EIDLE), 
        .PHY_REFCLK_MODE             (PHY_REFCLK_MODE),
        .PHY_REFCLK_FREQ             (PHY_REFCLK_FREQ)
    )
    cdr_ctrl_on_eidle_smsw_i
    (
        //----------------------------------------------------------------------------
        //  Input Ports
        //----------------------------------------------------------------------------
        .CDRCTRL_PCLK                               (pclk2_gt),
        .CDRCTRL_PCLK_RST_N                         (rst_psrst_n_r[3]),
        .CDRCTRL_CLK                                (PHY_REFCLK),
        .CDRCTRL_RST_N                              (rst_idle),
        .CDRCTRL_RATE                               (PHY_RATE),
        .CDRCTRL_RXELECIDLE                         (gt_rxelecidle[i]),
        .CDRCTRL_GEN34_EIOS_DET                     (gt_gen34_eios_det[i]),
        .CDRCTRL_RXCDRHOLD_IN                       (PHY_RXCDRHOLD),
        .CDRCTRL_RXCDRFREQRESET_IN                  (1'b0),
        .CDRCTRL_RXRATEDONE                         (gt_rxratedone[i]),
        //----------------------------------------------------------------------------
        //  Output Ports
        //----------------------------------------------------------------------------  
        .CDRCTRL_RXCDRHOLD_OUT                      (cdrctrl_rxcdrhold[i]),
        .CDRCTRL_RXCDRFREQRESET_OUT                 (cdrctrl_rxcdrfreqreset[i]),
        .CDRCTRL_RESETOVRD_OUT                      (cdrctrl_resetovrd[i])
    );
      
    assign gt_rxcdrhold[i] = (PHY_GEN12_CDR_CTRL_ON_EIDLE == "TRUE") || (PHY_GEN34_CDR_CTRL_ON_EIDLE == "TRUE") ? cdrctrl_rxcdrhold[i] : PHY_RXCDRHOLD;
    
    //----------------------------------------------------------------------------------------------
    //  Use Static GT Wrapper
    //----------------------------------------------------------------------------------------------
    if (PHY_GTWIZARD == "FALSE")
    
        begin : gt_wrapper_smsw
    
        //----------------------------------------------------------------------
        //  GT Channel
        //----------------------------------------------------------------------
        xp4_usp_smsw_gt_gt_channel #
        (
            .PHY_SIM_EN                     (PHY_SIM_EN),   
            .PHY_GT_XCVR                    (PHY_GT_XCVR),
            .PHY_MODE                       (PHY_MODE),
            .PHY_REFCLK_MODE                (PHY_REFCLK_MODE),
            .PHY_LANE                       (PHY_LANE),    
            .PHY_MAX_SPEED                  (PHY_MAX_SPEED),
            .PHY_GEN4_64BIT_EN              (PHY_GEN4_64BIT_EN),
            .PHY_GEN12_CDR_CTRL_ON_EIDLE     (PHY_GEN12_CDR_CTRL_ON_EIDLE),
            .PHY_GEN34_CDR_CTRL_ON_EIDLE     (PHY_GEN34_CDR_CTRL_ON_EIDLE),
            .PHY_REFCLK_FREQ                (PHY_REFCLK_FREQ),    
            .PHY_CORECLK_FREQ               (PHY_CORECLK_FREQ),         
            .GT_LANE_NUM                    (i)                      
        )
        gt_channel_smsw_i
        (  
        
            //------------------------------------------------------------------
            //  Clock Ports
            //------------------------------------------------------------------
            .GT_GTREFCLK0                   (PHY_GTREFCLK),
            .GT_TXUSRCLK                    (pclk),
            .GT_RXUSRCLK                    (pclk), 
            .GT_TXUSRCLK2                   (pclk2_gt),
            .GT_RXUSRCLK2                   (pclk2_gt), 
            
            .GT_TXOUTCLK                    (gt_txoutclk[i]), 
            .GT_RXOUTCLK                    (DBG_RXOUTCLK[i]), 
            .GT_TXOUTCLKFABRIC              (DBG_TXOUTCLKFABRIC[i]),                                                        
            .GT_RXOUTCLKFABRIC              (DBG_RXOUTCLKFABRIC[i]),                                                        
            .GT_TXOUTCLKPCS                 (DBG_TXOUTCLKPCS[i]),                                                        
            .GT_RXOUTCLKPCS                 (DBG_RXOUTCLKPCS[i]),  
            .GT_RXRECCLKOUT                 (DBG_RXRECCLKOUT[i]),
            
	    .GT_TXOUTCLKSEL                 (PHY_TXOUTCLKSEL),

            //------------------------------------------------------------------
            //  BUFG_GT Controller Ports                                               
            //------------------------------------------------------------------ 
            .GT_BUFGTCE                     (gt_bufgtce[i]),     
            .GT_BUFGTCEMASK                 (gt_bufgtcemask[(3*i)+2:(3*i)]), 
            .GT_BUFGTRESET                  (gt_bufgtreset[i]),
            .GT_BUFGTRSTMASK                (gt_bufgtrstmask[(3*i)+2:(3*i)]),   
            .GT_BUFGTDIV                    (gt_bufgtdiv[(9*i)+8:(9*i)]),
            
            //------------------------------------------------------------------
            //  Reset Ports
            //------------------------------------------------------------------
            .GT_CPLLPD                      (rst_cpllpd),
            .GT_CPLLRESET                   (rst_cpllreset),
            .GT_TXPROGDIVRESET              (rst_txprogdivreset),
            .GT_GTTXRESET                   (rst_gtreset),
            .GT_GTRXRESET                   (rst_gtreset), 
            .GT_TXUSERRDY                   (rst_userrdy),
            .GT_RXUSERRDY                   (rst_userrdy),              
                             
            .GT_TXPMARESET                  (DBG_TXPMARESET[i]),                                            
            .GT_RXPMARESET                  (DBG_RXPMARESET[i]),                                            
            .GT_TXPCSRESET                  (DBG_TXPCSRESET[i]),   
            .GT_RXPCSRESET                  (DBG_RXPCSRESET[i]),  
            .GT_RXBUFRESET                  (DBG_RXBUFRESET[i]),
            .GT_RXCDRRESET                  (DBG_RXCDRRESET[i]),  
            .GT_RXDFELPMRESET               (DBG_RXDFELPMRESET[i]), 
            .GT_RXCDRFREQRESET              (cdrctrl_rxcdrfreqreset[i]),
            
            .GT_RESETOVRD                   (cdrctrl_resetovrd[i]),
                             
            .GT_GTPOWERGOOD                 (gt_gtpowergood[i]), 
            .GT_TXPROGDIVRESETDONE          (gt_txprogdivresetdone[i]),     
            .GT_TXPMARESETDONE              (DBG_TXPMARESETDONE[i]),     
            .GT_RXPMARESETDONE              (DBG_RXPMARESETDONE[i]),             
            .GT_TXRESETDONE                 (gt_txresetdone[i]),
            .GT_RXRESETDONE                 (gt_rxresetdone[i]),                

            //------------------------------------------------------------------
            //  QPLL Ports
            //------------------------------------------------------------------
            .GT_QPLL0CLK                    (gtcom_qpll0outclk[i>>2]),                       
            .GT_QPLL0REFCLK                 (gtcom_qpll0outrefclk[i>>2]), 
            .GT_QPLL0LOCK                   (qpll0lock_all),                    // From all lanes
            .GT_QPLL1CLK                    (gtcom_qpll1outclk[i>>2]),
            .GT_QPLL1REFCLK                 (gtcom_qpll1outrefclk[i>>2]), 
            .GT_QPLL1LOCK                   (qpll1lock_all),                    // From all lanes
            
            .GT_QPLLRATE                    (gt_qpllrate[(3*i)+2:(3*i)]),
            
            //------------------------------------------------------------------
            //  Serial Line Ports
            //------------------------------------------------------------------
            .GT_RXP                         (PHY_RXP[i]),
            .GT_RXN                         (PHY_RXN[i]),
            
            .GT_TXP                         (PHY_TXP[i]),
            .GT_TXN                         (PHY_TXN[i]),
            
            //------------------------------------------------------------------
            //  TX Data Ports
            //------------------------------------------------------------------
            .GT_TXDATA                      (PHY_TXDATA[(64*i)+63:(64*i)]),
            .GT_TXDATAK                     (PHY_TXDATAK[(2*i)+1:(2*i)]),
            .GT_TXDATA_VALID                (PHY_TXDATA_VALID[i]),
            .GT_TXSTART_BLOCK               (PHY_TXSTART_BLOCK[i]),
            .GT_TXSYNC_HEADER               (PHY_TXSYNC_HEADER[(2*i)+1:(2*i)]),
            
            //------------------------------------------------------------------
            //  RX Data Ports
            //------------------------------------------------------------------
            .GT_RXDATA                      (PHY_RXDATA[(64*i)+63:(64*i)]),
            .GT_RXDATAK                     (PHY_RXDATAK[(2*i)+1:(2*i)]),
            .GT_RXDATA_VALID                (PHY_RXDATA_VALID[i]),
            .GT_RXSTART_BLOCK               (PHY_RXSTART_BLOCK[(2*i)+1:(2*i)]),
            .GT_RXSYNC_HEADER               (PHY_RXSYNC_HEADER[(2*i)+1:(2*i)]),
            
            //------------------------------------------------------------------
            //  PHY Command Ports
            //------------------------------------------------------------------
            .GT_TXDETECTRX                  (PHY_TXDETECTRX),
            .GT_TXELECIDLE                  (PHY_TXELECIDLE[i]), 
            .GT_TXCOMPLIANCE                (PHY_TXCOMPLIANCE[i]),
            .GT_RXPOLARITY                  (PHY_RXPOLARITY[i]),
            .GT_POWERDOWN                   (PHY_POWERDOWN),
            .GT_RATE                        (PHY_RATE), 
            .GT_RXCDRHOLD                   (gt_rxcdrhold[i]),      
                
            //------------------------------------------------------------------
            //  PHY Status Ports
            //------------------------------------------------------------------
            .GT_RXVALID                     (PHY_RXVALID[i]),
            .GT_PHYSTATUS                   (gt_phystatus[i]),
            .GT_RXELECIDLE                  (gt_rxelecidle[i]),
            .GT_RXSTATUS                    (PHY_RXSTATUS[(3*i)+2:(3*i)]),
                
            //------------------------------------------------------------------
            //  TX Driver Ports
            //------------------------------------------------------------------
            .GT_TXMARGIN                    (PHY_TXMARGIN),
            .GT_TXSWING                     (PHY_TXSWING),
            .GT_TXDEEMPH                    (PHY_TXDEEMPH),  
            
            //------------------------------------------------------------------
            //  TX Equalization Ports (Gen3) 
            //------------------------------------------------------------------
            .GT_TXPRECURSOR                 (txeq_precursor[(5*i)+4:(5*i)]),
            .GT_TXMAINCURSOR                (txeq_maincursor[(7*i)+6:(7*i)]),
            .GT_TXPOSTCURSOR                (txeq_postcursor[(5*i)+4:(5*i)]),
            
            //------------------------------------------------------------------
            //  PCIe Ports (Advance feature)
            //------------------------------------------------------------------
            .GT_PCIERSTIDLE                 (rst_idle),        
            .GT_PCIERSTTXSYNCSTART          (rst_txsync_start), 
            .GT_PCIEEQRXEQADAPTDONE         (1'd0),                             // Not used in top level
            .GT_PCIEUSERRATEDONE            (DBG_RATE_DONE[i]),                 // For debug only
        
            .GT_PCIEUSERPHYSTATUSRST        (gt_pcieuserphystatusrst[i]),    
            .GT_PCIERATEQPLLPD              (gt_pcierateqpllpd[(2*i)+1:(2*i)]),     
            .GT_PCIERATEQPLLRESET           (gt_pcierateqpllreset[(2*i)+1:(2*i)]), 
            .GT_PCIERATEIDLE                (gt_pcierateidle[i]),            
            .GT_PCIESYNCTXSYNCDONE          (gt_pciesynctxsyncdone[i]),  
            .GT_PCIERATEGEN3                (gt_pcierategen3[i]),               // Not used in top level
            .GT_PCIEUSERGEN3RDY             (gt_pcieusergen3rdy[i]),            // Not used in top level
            .GT_PCIEUSERRATESTART           (gt_pcieuserratestart[i]),          // For debug
            
            //------------------------------------------------------------------
            //  USB Ports
            //------------------------------------------------------------------
            .GT_TXONESZEROS                 (USB_TXONESZEROS[i]),                        
            .GT_RXEQTRAINING                (USB_RXEQTRAINING[i]),                       
            .GT_RXTERMINATION               (gt_rxtermination[i]),                        
    
            .GT_POWERPRESENT                (USB_POWERPRESENT[i]),    
            
            //------------------------------------------------------------------
            //  TX Sync Alignment Ports
            //------------------------------------------------------------------
            .GT_TXSYNCALLIN                 (txsyncallin_all),                  // From all lanes
            .GT_TXSYNCIN                    (gt_txsyncout[0]),                  // From master lane 0        
        
            .GT_TXPHALIGNDONE               (gt_txphaligndone[i]),            
            .GT_TXSYNCOUT                   (gt_txsyncout[i]),
            
             //-----------------------------------------------------------------
             //  Loopback and PRBS Ports
             //-----------------------------------------------------------------  
            .GT_LOOPBACK                    (DBG_LOOPBACK),                                              
            .GT_PRBSSEL                     (DBG_PRBSSEL),
            .GT_TXPRBSFORCEERR              (DBG_TXPRBSFORCEERR), 
            .GT_RXPRBSCNTRESET              (DBG_RXPRBSCNTRESET),                                                                                                      
        
            .GT_RXPRBSERR                   (DBG_RXPRBSERR[i]),                                              
            .GT_RXPRBSLOCKED                (DBG_RXPRBSLOCKED[i]),  
        
            //------------------------------------------------------------------
            //  GT Status Ports
            //------------------------------------------------------------------                                              
            .GT_MASTER_CPLLLOCK             (gt_cplllock[0]),                   // From master lane 0 
            
            .GT_CPLLLOCK                    (gt_cplllock[i]),  
            .GT_RXCDRLOCK                   (gt_rxcdrlock[i]),
            .GT_GEN34_EIOS_DET              (gt_gen34_eios_det[i]),
            .GT_RXRATEDONE                  (gt_rxratedone[i]),
            
            //------------------------------------------------------------------
            //  DRP Ports
            //------------------------------------------------------------------
            .GT_DRPCLK                      (PHY_REFCLK),
            .GT_DRPADDR                     (10'd0),
            .GT_DRPEN                       (1'b0),
            .GT_DRPWE                       (1'b0),
            .GT_DRPDI                       (16'd0),

            .GT_DRPRDY                      (),
            .GT_DRPDO                       ()            
        );
end // gt_channel            
        //------------------------------------------------------------------------------------------
        //  PHY Quad - Generate one Quad for every four Lanes
        //------------------------------------------------------------------------------------------
        if ((i%4)==0) 
                       
            begin : phy_quad   
                 
            //------------------------------------------------------------------
            //  Generate QPLL Powerdown and Reset
            //------------------------------------------------------------------
            //  * QPLL reset and powerdown for Quad 1 driven by       Master Lane 0
            //  * QPLL reset and powerdown for Quad 2 driven by Local Master Lane 4
            //------------------------------------------------------------------        
            assign qpll1pd[i>>2]    = (PHY_MAX_SPEED != 3) ? 1'd1 : (i > 3) ? (rst_qpllpd    || gt_pcierateqpllpd[(i*2)+1]) : 
                                                                              (rst_qpllpd    || gt_pcierateqpllpd[1]);
                                             
            assign qpll1reset[i>>2] = (PHY_MAX_SPEED != 3) ? 1'd1 : (i > 3) ? (rst_qpllreset || gt_pcierateqpllreset[(i*2)+1]) : 
                                                                              (rst_qpllreset || gt_pcierateqpllreset[1]);            
            
            assign qpll0pd[i>>2]    = (PHY_MAX_SPEED != 4) ? 1'd1 : (i > 3) ? (rst_qpllpd    || gt_pcierateqpllpd[(i*2)+0]) : 
                                                                              (rst_qpllpd    || gt_pcierateqpllpd[0]);
                                             
            assign qpll0reset[i>>2] = (PHY_MAX_SPEED != 4) ? 1'd1 : (i > 3) ? (rst_qpllreset || gt_pcierateqpllreset[(i*2)+0]) : 
                                                                              (rst_qpllreset || gt_pcierateqpllreset[0]);                                 
        
    if (PHY_GTWIZARD == "FALSE") begin : gt_common_smsw_int
            //------------------------------------------------------------------
            //  GT Common Module                                                   
            //------------------------------------------------------------------
            xp4_usp_smsw_gt_gt_common #
            (
                //--------------------------------------------------------------
                //  User Attributes
                //--------------------------------------------------------------
                .PHY_SIM_EN                 (PHY_SIM_EN),   
                .PHY_GT_XCVR                (PHY_GT_XCVR),
                .PHY_MAX_SPEED              (PHY_MAX_SPEED),
                .PHY_REFCLK_FREQ            (PHY_REFCLK_FREQ)          
            )
            gt_common_smsw_i
            (    
                //--------------------------------------------------------------
                //  Clock Ports
                //--------------------------------------------------------------
                .GTCOM_REFCLK               (PHY_GTREFCLK),
                
                .GTCOM_QPLL0LOCK            (gtcom_qpll0lock[i>>2]),
                .GTCOM_QPLL0OUTCLK          (gtcom_qpll0outclk[i>>2]),
                .GTCOM_QPLL0OUTREFCLK       (gtcom_qpll0outrefclk[i>>2]),
                
                .GTCOM_QPLL1LOCK            (gtcom_qpll1lock[i>>2]),
                .GTCOM_QPLL1OUTCLK          (gtcom_qpll1outclk[i>>2]),
                .GTCOM_QPLL1OUTREFCLK       (gtcom_qpll1outrefclk[i>>2]),
                
                //--------------------------------------------------------------
                //  Reset Ports
                //--------------------------------------------------------------             
                .GTCOM_QPLL0PD              (qpll0pd[i>>2]),         
                .GTCOM_QPLL0RESET           (qpll0reset[i>>2]),
                
                .GTCOM_QPLL1PD              (qpll1pd[i>>2]),         
                .GTCOM_QPLL1RESET           (qpll1reset[i>>2]),
                
                //--------------------------------------------------------------
                //  PCIe Ports
                //--------------------------------------------------------------    
                .GTCOM_QPLLRATE             ({1'd0, PHY_RATE}),               
                
                //--------------------------------------------------------------
                //  DRP Ports
                //--------------------------------------------------------------
                .GTCOM_DRPCLK               (GT_DRPCLK),                                     
                .GTCOM_DRPADDR              (GTCOM_DRPADDR[(16*(i>>2))+15:(16*(i>>2))]),                        
                .GTCOM_DRPEN                (GTCOM_DRPEN[i>>2]),                             
                .GTCOM_DRPWE                (GTCOM_DRPWE[i>>2]),
                .GTCOM_DRPDI                (GTCOM_DRPDI[(16*(i>>2))+15:(16*(i>>2))]),                     
                                                                             
                .GTCOM_DRPRDY               (GTCOM_DRPRDY[i>>2]),
                .GTCOM_DRPDO                (GTCOM_DRPDO[(16*(i>>2))+15:(16*(i>>2))])
            );
           end // gt_common_int

            end // phy_quad 
            
        end // phy_lane
       
endgenerate 
//--------------------------------------------------------------------------------------------------
//  Generate - End
//--------------------------------------------------------------------------------------------------
generate
    if (PHY_GTWIZARD == "TRUE") begin :gt_wizard_smsw

xp4_usp_smsw_gtwizard_top #
        (
            .PHY_LANE                       (PHY_LANE),                    
            .PHY_MAX_SPEED                  (PHY_MAX_SPEED),
            .PHY_GT_XCVR                    (PHY_GT_XCVR)
        )
        gtwizard_top_smsw_i
        (  
        
            //------------------------------------------------------------------
            //  Clock Ports *
            //------------------------------------------------------------------
            .GT_GTREFCLK0                   (PHY_GTREFCLK),                     
            .GT_TXUSRCLK                    ({PHY_LANE{pclk}}),
            .GT_RXUSRCLK                    ({PHY_LANE{pclk}}), 
            .GT_TXUSRCLK2                   ({PHY_LANE{pclk2_gt}}),
            .GT_RXUSRCLK2                   ({PHY_LANE{pclk2_gt}}), 
            
            .GT_RXOUTCLK                    (DBG_RXOUTCLK), 
            .GT_TXOUTCLKFABRIC              (DBG_TXOUTCLKFABRIC),                                                        
            .GT_RXOUTCLKFABRIC              (DBG_RXOUTCLKFABRIC),                                                        
            .GT_TXOUTCLKPCS                 (DBG_TXOUTCLKPCS),                                                        
            .GT_RXOUTCLKPCS                 (DBG_RXOUTCLKPCS),  
            .GT_RXRECCLKOUT                 (DBG_RXRECCLKOUT),
            .GT_TXOUTCLKSEL                 ({PHY_LANE{PHY_TXOUTCLKSEL}}),
            //------------------------------------------------------------------
            //  BUFG_GT Controller Ports *                                               
            //------------------------------------------------------------------ 
            .GT_BUFGTCE                     (gt_bufgtce),     
            .GT_BUFGTCEMASK                 (gt_bufgtcemask), 
            .GT_BUFGTRESET                  (gt_bufgtreset),
            .GT_BUFGTRSTMASK                (gt_bufgtrstmask),   
            .GT_BUFGTDIV                    (gt_bufgtdiv),
            .GT_TXOUTCLK                    (gt_txoutclk),   
            
            //------------------------------------------------------------------  
            //  Reset Ports *                                                      
            //------------------------------------------------------------------  
            .GT_CPLLPD                      ({PHY_LANE{rst_cpllpd}}),              
            .GT_CPLLRESET                   ({PHY_LANE{rst_cpllreset}}),           
            .GT_TXPROGDIVRESET              ({PHY_LANE{rst_txprogdivreset}}),        
            .GT_RXPROGDIVRESET              ({PHY_LANE{rst_txprogdivreset}}),        
            .GT_GTTXRESET                   ({PHY_LANE{rst_gtreset}}),             
            .GT_GTRXRESET                   ({PHY_LANE{rst_gtreset}}),             
            .GT_TXUSERRDY                   ({PHY_LANE{rst_userrdy}}),             
            .GT_RXUSERRDY                   ({PHY_LANE{rst_userrdy}}),             
                                                                                  
            .GT_TXPMARESET                  (DBG_TXPMARESET),                                            
            .GT_RXPMARESET                  (DBG_RXPMARESET),                                            
            .GT_TXPCSRESET                  (DBG_TXPCSRESET),   
            .GT_RXPCSRESET                  (DBG_RXPCSRESET),  
            .GT_RXBUFRESET                  (DBG_RXBUFRESET),
            .GT_RXCDRRESET                  (DBG_RXCDRRESET),  
            .GT_RXDFELPMRESET               (DBG_RXDFELPMRESET),                                

            .GT_GTPOWERGOOD                 (gt_gtpowergood),                     
            .GT_TXPROGDIVRESETDONE          (gt_txprogdivresetdone),              
            .GT_TXRESETDONE                 (gt_txresetdone),                     
            .GT_RXRESETDONE                 (gt_rxresetdone),                     
            .GT_TXPMARESETDONE              (DBG_TXPMARESETDONE),     
            .GT_RXPMARESETDONE              (DBG_RXPMARESETDONE),             
            
            //--------------------------------------------------------------
            //  Common QPLL Ports *
            //--------------------------------------------------------------
            .GTCOM_QPLLPD                   (rst_qpllpd),         
            .GTCOM_QPLLRESET                (rst_qpllreset), 
            
            .GTCOM_QPLL1LOCK                (gtcom_qpll1lock),
            .GTCOM_QPLL0LOCK                (gtcom_qpll0lock),

            .GTCOM_QPLL0OUTCLK              (gtcom_qpll0outclk),
            .GTCOM_QPLL0OUTREFCLK           (gtcom_qpll0outrefclk),
            .GTCOM_QPLL1OUTCLK              (gtcom_qpll1outclk),
            .GTCOM_QPLL1OUTREFCLK           (gtcom_qpll1outrefclk),
            //--------------------------------------------------------------
            //  Common DRP Ports *
            //--------------------------------------------------------------
            .GTCOM_DRPCLK                   (GT_DRPCLK),                                     
            .GTCOM_DRPADDR                  (GTCOM_DRPADDR),                        
            .GTCOM_DRPEN                    (GTCOM_DRPEN),                             
            .GTCOM_DRPWE                    (GTCOM_DRPWE),
            .GTCOM_DRPDI                    (GTCOM_DRPDI),                     
                                                                             
            .GTCOM_DRPRDY                   (GTCOM_DRPRDY),
            .GTCOM_DRPDO                    (GTCOM_DRPDO),

            .GT_DRPCLK                      ({PHY_LANE{PHY_REFCLK}}),
            .GT_DRPADDR                     (gt_drpaddr),
            .GT_DRPEN                       (gt_drpen),
            .GT_DRPWE                       (gt_drpwe),
            .GT_DRPDI                       (gt_drpdi),

            .GT_DRPRDY                      (gt_drprdy),
            .GT_DRPDO                       (gt_drpdo),            
            //------------------------------------------------------------------
            //  Serial Line Ports *
            //------------------------------------------------------------------
            .GT_RXP                         (PHY_RXP),
            .GT_RXN                         (PHY_RXN),
            
            .GT_TXP                         (PHY_TXP),
            .GT_TXN                         (PHY_TXN),
            
            //------------------------------------------------------------------
            //  TX Data Ports *
            //------------------------------------------------------------------
            .GT_TXDATA                      (PHY_TXDATA),
            .GT_TXDATAK                     (PHY_TXDATAK),
            .GT_TXDATA_VALID                (PHY_TXDATA_VALID),
            .GT_TXSTART_BLOCK               (PHY_TXSTART_BLOCK),
            .GT_TXSYNC_HEADER               (PHY_TXSYNC_HEADER),
            
            //------------------------------------------------------------------
            //  RX Data Ports *
            //------------------------------------------------------------------
            .GT_RXDATA                      (PHY_RXDATA),
            .GT_RXDATAK                     (PHY_RXDATAK),
            .GT_RXDATA_VALID                (PHY_RXDATA_VALID),
            .GT_RXSTART_BLOCK               (PHY_RXSTART_BLOCK),
            .GT_RXSYNC_HEADER               (PHY_RXSYNC_HEADER),
            
            //------------------------------------------------------------------
            //  PHY Command Ports *
            //------------------------------------------------------------------
            .GT_TXDETECTRX                  ({PHY_LANE{PHY_TXDETECTRX}}),
            .GT_TXELECIDLE                  (PHY_TXELECIDLE), 
            .GT_TXCOMPLIANCE                (PHY_TXCOMPLIANCE),
            .GT_RXPOLARITY                  (PHY_RXPOLARITY),
            .GT_POWERDOWN                   ({PHY_LANE{PHY_POWERDOWN}}),
            .GT_RATE                        ({PHY_LANE{PHY_RATE}}),       
            .GT_RXCDRHOLD                   (gt_rxcdrhold),      
                
            //------------------------------------------------------------------
            //  PHY Status Ports *
            //------------------------------------------------------------------
            .GT_RXVALID                     (PHY_RXVALID),
            .GT_PHYSTATUS                   (gt_phystatus),
            .GT_RXELECIDLE                  (gt_rxelecidle),
            .GT_RXSTATUS                    (PHY_RXSTATUS),
                
            //------------------------------------------------------------------
            //  TX Driver Ports *
            //------------------------------------------------------------------
            .GT_TXMARGIN                    ({PHY_LANE{PHY_TXMARGIN}}),
            .GT_TXSWING                     ({PHY_LANE{PHY_TXSWING}}),
            .GT_TXDEEMPH                    ({PHY_LANE{PHY_TXDEEMPH}}),  
            
            //------------------------------------------------------------------
            //  TX Equalization Ports (Gen3) *
            //------------------------------------------------------------------
            .GT_TXPRECURSOR                 (txeq_precursor),
            .GT_TXMAINCURSOR                (txeq_maincursor),
            .GT_TXPOSTCURSOR                (txeq_postcursor),
            
            //------------------------------------------------------------------
            //  PCIe PCS (Advance Feature) *
            //------------------------------------------------------------------
            .GT_PCIERSTIDLE                 ({PHY_LANE{rst_idle}}),        
            .GT_PCIERSTTXSYNCSTART          ({PHY_LANE{rst_txsync_start}}), 
            .GT_PCIEEQRXEQADAPTDONE         ({PHY_LANE{1'd0}}),                 // Not used
            .GT_PCIEUSERRATEDONE            (DBG_RATE_DONE),                 // For debug only
        
            .GT_PCIEUSERPHYSTATUSRST        (gt_pcieuserphystatusrst),    
            .GT_PCIERATEQPLLPD              (gt_pcierateqpllpd),     
            .GT_PCIERATEQPLLRESET           (gt_pcierateqpllreset), 
            .GT_PCIERATEIDLE                (gt_pcierateidle),            
            .GT_PCIESYNCTXSYNCDONE          (gt_pciesynctxsyncdone),  
            .GT_PCIERATEGEN3                (gt_pcierategen3),    
            .GT_PCIEUSERGEN3RDY             (gt_pcieusergen3rdy),  
            .GT_PCIEUSERRATESTART           (gt_pcieuserratestart), 
            
            .GT_TXPHALIGNDONE               (gt_txphaligndone),            
             //-----------------------------------------------------------------
             //  Loopback and PRBS Ports *
             //-----------------------------------------------------------------  
						.GT_LOOPBACK                    ({PHY_LANE{DBG_LOOPBACK}}),                                              
            .GT_PRBSSEL                     ({PHY_LANE{DBG_PRBSSEL}}),
            .GT_TXPRBSFORCEERR              ({PHY_LANE{DBG_TXPRBSFORCEERR}}), 
            .GT_TXINHIBIT                   ({PHY_LANE{1'd0}}),
            .GT_RXPRBSCNTRESET              ({PHY_LANE{DBG_RXPRBSCNTRESET}}),                                                                                                      
            
            .GT_RXPRBSERR                   (DBG_RXPRBSERR),                                              
            .GT_RXPRBSLOCKED                (DBG_RXPRBSLOCKED),  
        
            .GT_TXDLYSRESETDONE             ( ),//(GT_TXDLYSRESETDONE ),    
            .GT_TXPHINITDONE                ( ),//(GT_TXPHINITDONE),
            .GT_RXCOMMADET                  ( ),//(GT_RXCOMMADET),
            .GT_RXBUFSTATUS                 ( ),//(GT_RXBUFSTATUS),
            //------------------------------------------------------------------
            //  GT Status Ports *
            //------------------------------------------------------------------                                                   
            .GT_CPLLLOCK                    (gt_cplllock),  
            .GT_RXCDRLOCK                   (gt_rxcdrlock),

            .GT_GEN34_EIOS_DET              (gt_gen34_eios_det),
            .GT_RXRATEDONE                  (gt_rxratedone),

            //------------------------------------------------------------------
            //  GT RX Termination
            //------------------------------------------------------------------   
            .GT_RXTERMINATION               (gt_rxtermination)
        );
    end
endgenerate 

//--------------------------------------------------------------------------------------------------
//  Convert per-lane signals to per-design 
//--------------------------------------------------------------------------------------------------
    assign qpll0lock_all   = &gtcom_qpll0lock;
    assign qpll1lock_all   = &gtcom_qpll1lock;
    assign txsyncallin_all = &gt_txphaligndone;

//------------------------------------------------------------------------------
//  PHYSTATUS Reset Synchronizer for PCLK 
//------------------------------------------------------------------------------

always @ (posedge pclk or negedge rst_idle)
  begin
    if (!rst_idle)
      rst_psrst_n_r <= 4'd0;
    else
      rst_psrst_n_r <= {rst_psrst_n_r[2:0], 1'd1};
  end

//--------------------------------------------------------------------------------------------------
//  PHY Wrapper Outputs
//--------------------------------------------------------------------------------------------------
assign PHY_PCLK               = pclk;
assign PHY_PHYSTATUS          = gt_phystatus;
assign PHY_PHYSTATUS_RST      = !rst_psrst_n_r[3];
assign PHY_RXELECIDLE         = gt_rxelecidle;

//------------------------------------------------------------------------------
//  TX Equalization Outputs (Gen3/Gen4) 
//------------------------------------------------------------------------------
assign PHY_TXEQ_FS            = 6'd40;                                          // Value based on GT TX driver characteristic                                    
assign PHY_TXEQ_LF            = 6'd12;                                          // Value based on GT TX driver characteristic
assign PHY_TXEQ_NEW_COEFF     = txeq_new_coeff;        
assign PHY_TXEQ_DONE          = txeq_done;                                                   
      
//------------------------------------------------------------------------------
//  RX Equalization Outputs (Gen3/Gen4)
//------------------------------------------------------------------------------     
assign PHY_RXEQ_LFFS_SEL      = rxeq_lffs_sel;                                                  
assign PHY_RXEQ_NEW_TXCOEFF   = rxeq_new_txcoeff;     
assign PHY_RXEQ_ADAPT_DONE    = rxeq_adapt_done;   
assign PHY_RXEQ_DONE          = rxeq_done;   

//------------------------------------------------------------------------------
//  Debug Outputs 
//------------------------------------------------------------------------------ 
assign DBG_RATE_START         = gt_pcieuserratestart;
assign DBG_RST_IDLE           = rst_idle;
assign DBG_RATE_IDLE          = gt_pcierateidle;
assign DBG_RXCDRLOCK          = gt_rxcdrlock;     

assign DBG_TXOUTCLK           = gt_txoutclk;     
    
assign DBG_RRST_N             = rrst_n;
assign DBG_PRST_N             = prst_n;
assign DBG_GTPOWERGOOD        = gt_gtpowergood;
assign DBG_CPLLLOCK           = gt_cplllock;
assign DBG_QPLL0LOCK          = gtcom_qpll0lock;
assign DBG_QPLL1LOCK          = gtcom_qpll1lock;
assign DBG_TXPROGDIVRESETDONE = gt_txprogdivresetdone;
assign DBG_TXRESETDONE        = gt_txresetdone;
assign DBG_RXRESETDONE        = gt_rxresetdone;
assign DBG_TXSYNCDONE         = gt_pciesynctxsyncdone;
assign DBG_GEN34_EIOS_DET     = gt_gen34_eios_det;
                                           
           

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_gt_cdr_ctrl_on_eidle.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
//  Design :  PHY Wrapper
//  Module :  CDR Control Upon EIDLE Detection
//--------------------------------------------------------------------------------------------------

`timescale 1ps / 1ps

//--------------------------------------------------------------------------------------------------
//  CDR Control Upon EIDLE Detection Module
//--------------------------------------------------------------------------------------------------
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_gt_cdr_ctrl_on_eidle #
(
    parameter         PHY_GEN12_CDR_CTRL_ON_EIDLE = "FALSE",
    parameter         PHY_GEN34_CDR_CTRL_ON_EIDLE = "FALSE",
    parameter integer PHY_REFCLK_MODE            = 0,
    parameter integer SYNC_STAGE                 = 3,
    parameter integer PHY_REFCLK_FREQ            = 0
)
(
    //-------------------------------------------------------------------------- 
    //  Input Ports
    //-------------------------------------------------------------------------- 
    input                               CDRCTRL_PCLK,
    input                               CDRCTRL_PCLK_RST_N,
    input                               CDRCTRL_CLK,
    input                               CDRCTRL_RST_N,
    input     [ 1:0]                    CDRCTRL_RATE,
    input                               CDRCTRL_RXELECIDLE,
    input                               CDRCTRL_GEN34_EIOS_DET,
    input                               CDRCTRL_RXCDRHOLD_IN,    
    input                               CDRCTRL_RXCDRFREQRESET_IN,
    input                               CDRCTRL_RXRATEDONE,
    
    //-------------------------------------------------------------------------- 
    //  Output Ports
    //-------------------------------------------------------------------------- 
    output                              CDRCTRL_RXCDRFREQRESET_OUT,
    output                              CDRCTRL_RXCDRHOLD_OUT,
    output                              CDRCTRL_RESETOVRD_OUT
);
    //--------------------------------------------------------------------------
    //  Synchronized Signals
    //--------------------------------------------------------------------------                                     
    wire                                gen3or4;
    reg         [ 1:0]                  rate_r;     
    reg         [ 1:0]                  rate_r2;
    wire                                rxelecidle_a;
    reg         [ 1:0]                  rxelecidle_r;
    wire                                gen34_eios_det_a;
    reg         [ 1:0]                  gen34_eios_det_r;
    wire                                rxcdrhold_in_r;
    reg                                 rate_change;
    wire                                rate_change_a;
    
    reg        [6:0]    rxelecidle_cycle_count;
    wire        ctrl_fsm_not_in_solid_deassert;
    //-------------------------------------------------------------------------- 
    //  FSM Signals
    //-------------------------------------------------------------------------- 
    reg [ 2:0] fsm;
    
    reg                                 rxcdrhold = 1'd0;     
    reg        [ 7:0]                   counter_max = 8'd0;
    reg        [ 7:0]                   wait_ctr = 8'd0;
    reg                                 resetovrd = 1'd0;
    reg                                 rxcdrfreqreset = 1'd0;
    
    reg                                 exit = 1'd0;
    wire                                rst_n;

    localparam MAX_COUNT_ENTER = (PHY_REFCLK_FREQ == 2) ? 8'd9 : 
                                 (PHY_REFCLK_FREQ == 1) ? 8'd4  : 8'd3;
    
    localparam MAX_COUNT_EXIT = (PHY_REFCLK_FREQ == 2)  ? 8'd75 : 
                                 (PHY_REFCLK_FREQ == 1) ? 8'd38 : 8'd30;
    
    assign rst_n = CDRCTRL_RST_N;

    reg [3:0] gen34_eios_det_extend;
    reg [7:0] rate_change_extend = 8'd0;
    reg rxelecidle_int = 0;
    reg gen34_eios_det_pclk;
    reg rate_change_extend_pclk;
    
    always @(posedge CDRCTRL_PCLK) 
    begin
      if (!CDRCTRL_PCLK_RST_N) begin
        gen34_eios_det_extend <= 4'd0;
        gen34_eios_det_pclk <= 1'd0;
      end 
      else begin
        gen34_eios_det_extend <= {gen34_eios_det_extend[2:0],CDRCTRL_GEN34_EIOS_DET};
        gen34_eios_det_pclk <= |gen34_eios_det_extend;
      end
    end
    
    //--------------------------------------------------------------------------------------------------
    //  Input Synchronizer or Pipeline
    //--------------------------------------------------------------------------------------------------
    xp4_usp_smsw_sync #(.WIDTH (1), .STAGE (SYNC_STAGE)) sync_gen34          (.CLK (CDRCTRL_CLK), .D (CDRCTRL_RATE[1]),         .Q (gen3or4));
    xp4_usp_smsw_sync #(.WIDTH (1), .STAGE (SYNC_STAGE)) sync_rxelecidle     (.CLK (CDRCTRL_CLK), .D (CDRCTRL_RXELECIDLE),      .Q (rxelecidle_a));
    xp4_usp_smsw_sync #(.WIDTH (1), .STAGE (SYNC_STAGE)) sync_gen34_eios_det (.CLK (CDRCTRL_CLK), .D (gen34_eios_det_pclk),     .Q (gen34_eios_det_a));
    xp4_usp_smsw_sync #(.WIDTH (1), .STAGE (SYNC_STAGE)) sync_rxcdrreset_in  (.CLK (CDRCTRL_CLK), .D (CDRCTRL_RXCDRHOLD_IN),    .Q (rxcdrhold_in_r));
    
    always @ (posedge CDRCTRL_CLK) 
    begin
      if (!rst_n) begin
        rxelecidle_r <= 2'd3;
        gen34_eios_det_r <= 2'd0;
      end 
      else begin 
        rxelecidle_r <= {rxelecidle_r[0], rxelecidle_a}; 
        gen34_eios_det_r <= {gen34_eios_det_r[0], gen34_eios_det_a}; 
      end
    end 
    
generate
    if (PHY_REFCLK_MODE <= 1) 
    begin : non_sris
    //--------------------------------------------------------------------------
    //  FSM Encoding
    //-------------------------------------------------------------------------- 
    localparam FSM_IDLE                  = 3'd0;
    localparam FSM_GEN12_RXELECIDLE_EXIT = 3'd1;
    localparam FSM_GEN34_RXELECIDLE_EXIT = 3'd2;

  assign ctrl_fsm_not_in_solid_deassert = (fsm == FSM_IDLE);
    
      always @ (posedge CDRCTRL_CLK) 
      begin 
        if (ctrl_fsm_not_in_solid_deassert) begin
          rxelecidle_cycle_count <= 7'd0;
        end 
        else begin
          if (!rxelecidle_r[1])
            rxelecidle_cycle_count <= rxelecidle_cycle_count + 7'd1;        
          else 
            rxelecidle_cycle_count <= 7'd0;
        end
      end
      
      always @(posedge CDRCTRL_CLK)
      begin 
        if (ctrl_fsm_not_in_solid_deassert) begin
          rxelecidle_int <= 1'b0;
        end 
        else begin
          if (rxelecidle_cycle_count > 64)
            rxelecidle_int <= 1'b1;
          else 
            rxelecidle_int <= rxelecidle_int;
        end
      end
    
    //--------------------------------------------------------------------------------------------------
    //  Hold CDR upon EIOS/EIDLE detection FSM
    //--------------------------------------------------------------------------------------------------
      always @ (posedge CDRCTRL_CLK)
      begin

          if (!rst_n)
              begin
              fsm        <= FSM_IDLE;
              rxcdrhold  <= 1'd0;
              end
          else
              begin
              
              case (fsm)
                  
              //------------------------------------------------------------------------------------------
              //  Stay in IDLE state until EIOS/EIDLE rising edge is detected
              //------------------------------------------------------------------------------------------
              FSM_IDLE :
              
                  begin
                 if ((PHY_GEN12_CDR_CTRL_ON_EIDLE == "TRUE") && (!gen3or4) && (!rxelecidle_r[1]&rxelecidle_r[0]))
                      begin
                      fsm       <= FSM_GEN12_RXELECIDLE_EXIT;
                      rxcdrhold <= 1'd1;
                      end
                 else if ((PHY_GEN34_CDR_CTRL_ON_EIDLE == "TRUE") && (gen3or4) && (!gen34_eios_det_r[1]&gen34_eios_det_r[0]))
                      begin
                      fsm       <= FSM_GEN34_RXELECIDLE_EXIT;
                      rxcdrhold <= 1'd1;
                      end
                  else
                      begin
                      fsm       <= FSM_IDLE;
                      rxcdrhold <= rxcdrhold_in_r;
                      end
                  end     
                  
              //------------------------------------------------------------------------------------------
              //  Gen1/Gen2:  Hold RXCDRRESET until RXELECIDLE exit
              //------------------------------------------------------------------------------------------
              FSM_GEN12_RXELECIDLE_EXIT:
              
                  begin
                  if (rxelecidle_int)
                      begin
                      fsm        <= FSM_IDLE;
                      rxcdrhold  <= 1'd0;
                      end
                  else
                      begin
                      fsm        <= FSM_GEN12_RXELECIDLE_EXIT;
                      rxcdrhold  <= 1'd1;
                      end
                  end    
                  
              //------------------------------------------------------------------------------------------
              //  Gen3/Gen4:  Hold RXCDRRESET until RXELECIDLE exit
              //------------------------------------------------------------------------------------------
              FSM_GEN34_RXELECIDLE_EXIT:
              
                  begin
                  if ((!gen34_eios_det_r[0]) & rxelecidle_int)
                      begin
                      fsm        <= FSM_IDLE;
                      rxcdrhold  <= 1'd0;
                      end
                  else
                      begin
                      fsm        <= FSM_GEN34_RXELECIDLE_EXIT;
                      rxcdrhold  <= 1'd1;
                      end
                  end    
                  
              //------------------------------------------------------------------------------------------
              //  Default State
              //------------------------------------------------------------------------------------------
              default :
              
                  begin
                  fsm        <= FSM_IDLE;
                  rxcdrhold <= 1'd0;
                  end

              endcase
              
              end
              
      end
    end 
endgenerate

generate
  if (PHY_REFCLK_MODE == 2) begin : sris
  
    reg [7:0]rx_rate_done_extend = 8'd0;
    reg rx_rate_done_extend_pclk = 1'd0;
    wire rate_done_a;
    reg rate_change_in_prog = 1'd0;
  
    always @(posedge CDRCTRL_PCLK)
    begin
      if (!CDRCTRL_PCLK_RST_N) begin
        rate_r <= 2'd0;
        rate_r2 <= 2'd0;
        rate_change <= 1'b0;
        rate_change_extend_pclk <= 1'd0;
        rate_change_extend <= 7'd0;
        rx_rate_done_extend_pclk <= 1'd0;
        rx_rate_done_extend <= 7'd0;        
      end
      else begin
        rate_r <= CDRCTRL_RATE;
        rate_r2 <= rate_r;

        if (rate_r2 != rate_r) 
          rate_change <= 1'b1;
        else
          rate_change <= 1'b0;
          
        rate_change_extend <= {rate_change_extend[6:0],rate_change};
        rate_change_extend_pclk <= |rate_change_extend;  

        rx_rate_done_extend <= {rx_rate_done_extend[6:0],CDRCTRL_RXRATEDONE};
        rx_rate_done_extend_pclk <= |rx_rate_done_extend;          
        
      end  
    end
    
    xp4_usp_smsw_sync #(.WIDTH (1), .STAGE (SYNC_STAGE)) sync_rate_change    (.CLK (CDRCTRL_CLK), .D (rate_change_extend_pclk), .Q (rate_change_a));
    xp4_usp_smsw_sync #(.WIDTH (1), .STAGE (SYNC_STAGE)) sync_rate_done      (.CLK (CDRCTRL_CLK), .D (rx_rate_done_extend_pclk), .Q (rate_done_a));
    
    //--------------------------------------------------------------------------
    //  FSM Encoding
    //-------------------------------------------------------------------------- 
    localparam FSM_IDLE                                 = 3'd0;
    localparam FSM_COUNTER                              = 3'd1;
    localparam FSM_GEN12_RXELECIDLE_EXIT_OR_RATE_CHANGE = 3'd2;
    localparam FSM_GEN34_RXELECIDLE_EXIT_OR_RATE_CHANGE = 3'd3;
    localparam FSM_WAIT_RATE_DONE                       = 3'd4;
    
    //--------------------------------------------------------------------------------------------------
    //  Reset CDR upon EIOS/EIDLE detection FSM
    //--------------------------------------------------------------------------------------------------
      always @ (posedge CDRCTRL_CLK)
      begin

          if (!rst_n)
              begin
              fsm            <= FSM_IDLE;
              resetovrd      <= 1'd0;
              rxcdrfreqreset <= 1'd0;
              wait_ctr       <= 8'd0;
              counter_max    <= 8'd0;
              exit           <= 1'd0;
              rate_change_in_prog <= 1'd0;
              end
          else
              begin
              
              case (fsm)
                  
              //------------------------------------------------------------------------------------------
              //  Stay in IDLE state until EIOS/EIDLE rising edge is detected
              //------------------------------------------------------------------------------------------
              FSM_IDLE :
              
                begin
                exit           <= 1'd0;
                
                counter_max <= MAX_COUNT_ENTER;
                
                 if ((PHY_GEN12_CDR_CTRL_ON_EIDLE == "TRUE") && ((!gen3or4) && (!rxelecidle_r[1]&rxelecidle_r[0])) || (rate_change_in_prog && !rxelecidle_r[0]) )
                      begin
                      fsm        <= FSM_COUNTER;
                      resetovrd  <= 1'd1;
                      rxcdrfreqreset <= 1'd0;
                      end
                 else if ((PHY_GEN34_CDR_CTRL_ON_EIDLE == "TRUE") && (gen3or4) && (!gen34_eios_det_r[1]&gen34_eios_det_r[0]) || (rate_change_in_prog && !rxelecidle_r[0]))
                      begin
                      fsm        <= FSM_COUNTER;
                      resetovrd  <= 1'd1;
                      rxcdrfreqreset <= 1'd0;
                      end
                  else
                      begin
                      fsm       <= FSM_IDLE;
                      resetovrd <= 1'd0;
                      rxcdrfreqreset <= 1'd0;
                      end
                      
                  end     
              
              FSM_COUNTER : 
              
                begin
                  if (wait_ctr < counter_max)
                  begin
                    wait_ctr <= wait_ctr + 1'b1;
                    fsm <= FSM_COUNTER;
                  end
                  else begin
                    wait_ctr <= 8'd0;
                    
                    if (!exit && !gen3or4) begin
                      rxcdrfreqreset <= 1'd1;
                      fsm <= FSM_GEN12_RXELECIDLE_EXIT_OR_RATE_CHANGE;
                    end
                    else if (!exit && gen3or4) begin
                      rxcdrfreqreset <= 1'd1;
                      fsm <= FSM_GEN34_RXELECIDLE_EXIT_OR_RATE_CHANGE;
                    end
                    else if (exit && rate_change_in_prog) begin
                      fsm <= FSM_WAIT_RATE_DONE;
                      resetovrd <= 1'd0;
                    end
                    else begin
                      fsm <= FSM_IDLE;
                      resetovrd <= 1'd0;
                    end
                  end
                end
              
              //------------------------------------------------------------------------------------------
              //  Gen1/Gen2:  Hold RXCDRREQRESET until RXELECIDLE exit or rate change detected
              //------------------------------------------------------------------------------------------
              FSM_GEN12_RXELECIDLE_EXIT_OR_RATE_CHANGE:
              
                  begin
                  
                  exit <= 1'd1;
                  
                  counter_max <= 8'd30;
                  
                  if (!rxelecidle_r[0] || rate_change_a)
                      begin
                      rate_change_in_prog <= rate_change_a;
                      fsm            <= FSM_COUNTER;
                      rxcdrfreqreset <= 1'd0;
                      end
                  else
                      begin
                      fsm        <= FSM_GEN12_RXELECIDLE_EXIT_OR_RATE_CHANGE;
                      end
                  end
                  
              //------------------------------------------------------------------------------------------
              //  Gen3/Gen4:  Hold RXCDRREQRESET until RXELECIDLE exit or rate change detected
              //------------------------------------------------------------------------------------------
              FSM_GEN34_RXELECIDLE_EXIT_OR_RATE_CHANGE:
                  begin 
 
                  exit <= 1'd1;
 
                  counter_max <= MAX_COUNT_EXIT;
                  
                  if (((!gen34_eios_det_r[0]) & (!rxelecidle_r[0])) || rate_change_a)
                      begin
                      rate_change_in_prog <= rate_change_a;
                      fsm            <= FSM_COUNTER;
                      rxcdrfreqreset <= 1'd0;
                      end
                  else
                      begin
                      fsm            <= FSM_GEN34_RXELECIDLE_EXIT_OR_RATE_CHANGE;
                      end
                  end    

              FSM_WAIT_RATE_DONE:
                begin 
                  
                  if (rate_done_a) 
                    fsm <= FSM_IDLE;
                  else 
                    fsm <= FSM_WAIT_RATE_DONE;
               
                end                  
              
              //------------------------------------------------------------------------------------------
              //  Default State
              //------------------------------------------------------------------------------------------
              default :
              
                  begin
                  fsm            <= FSM_IDLE;
                  resetovrd      <= 1'd0;
                  rxcdrfreqreset <= 1'd0;
                  wait_ctr       <= 8'd0;
                  counter_max    <= 8'd0;         
                  exit           <= 1'd0;
                  end

              endcase
              
              end
        end      
      end
endgenerate

//--------------------------------------------------------------------------------------------------
//  HOLD CDR upon EIOS/EIDLE Detection Outputs
//--------------------------------------------------------------------------------------------------
assign CDRCTRL_RXCDRHOLD_OUT = rxcdrhold;

//--------------------------------------------------------------------------------------------------
//  RESET CDR upon EIOS/EIDLE Detection Outputs
//--------------------------------------------------------------------------------------------------
assign CDRCTRL_RXCDRFREQRESET_OUT = rxcdrfreqreset;
assign CDRCTRL_RESETOVRD_OUT = resetovrd;


endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_gt_gt_channel.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
//  Design :  PHY Wrapper 
//  Module :  GT Channel
//--------------------------------------------------------------------------------------------------

`timescale 1ps / 1ps

//--------------------------------------------------------------------------------------------------
//  GT Channel Module
//--------------------------------------------------------------------------------------------------
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_gt_gt_channel #
(
    parameter         PHY_SIM_EN                 = "FALSE", 
    parameter         PHY_GT_XCVR                = "GTY",
    parameter integer PHY_MODE                   = 0,
    parameter integer PHY_REFCLK_MODE            = 0,
    parameter integer PHY_LANE                   = 1,
    parameter integer PHY_MAX_SPEED              = 3,
    parameter         PHY_GEN4_64BIT_EN          = "FALSE",
    parameter         PHY_GEN12_CDR_CTRL_ON_EIDLE = "FALSE",   
    parameter         PHY_GEN34_CDR_CTRL_ON_EIDLE = "FALSE", 
    parameter integer PHY_REFCLK_FREQ            = 0,                
    parameter integer PHY_CORECLK_FREQ           = 2,
    parameter         GT_LANE_NUM                = 0
)
(    
    //--------------------------------------------------------------------------
    //  Clock Ports
    //--------------------------------------------------------------------------
    input                               GT_GTREFCLK0,
    input                               GT_TXUSRCLK,
    input                               GT_RXUSRCLK,
    input                               GT_TXUSRCLK2,
    input                               GT_RXUSRCLK2,    

    output                              GT_TXOUTCLK, 
    output                              GT_RXOUTCLK,
    output                              GT_TXOUTCLKFABRIC,                                                        
    output                              GT_RXOUTCLKFABRIC,                                                        
    output                              GT_TXOUTCLKPCS,                                                        
    output                              GT_RXOUTCLKPCS,  
    output                              GT_RXRECCLKOUT,

    input       [ 2:0]                  GT_TXOUTCLKSEL,             
    
    //--------------------------------------------------------------------------   
    //  BUFG_GT Controller Ports                                                                        
    //--------------------------------------------------------------------------                   
    output                              GT_BUFGTCE,       
    output      [ 2:0]                  GT_BUFGTCEMASK, 
    output                              GT_BUFGTRESET,
    output      [ 2:0]                  GT_BUFGTRSTMASK,
    output      [ 8:0]                  GT_BUFGTDIV,   
                
    //--------------------------------------------------------------------------
    //  Reset Ports
    //--------------------------------------------------------------------------
    input                               GT_CPLLPD,
    input                               GT_CPLLRESET,
    input                               GT_TXPROGDIVRESET,
    input                               GT_GTTXRESET,
    input                               GT_GTRXRESET,
    input                               GT_TXUSERRDY,
    input                               GT_RXUSERRDY,
    
    input                               GT_TXPMARESET,                                            
    input                               GT_RXPMARESET,                                            
    input                               GT_TXPCSRESET,   
    input                               GT_RXPCSRESET,  
    input                               GT_RXBUFRESET,
    input                               GT_RXCDRRESET,
    input                               GT_RXDFELPMRESET,
    input                               GT_RXCDRFREQRESET,
    
    input                               GT_RESETOVRD,
                                        
    output                              GT_GTPOWERGOOD,
    output                              GT_TXPROGDIVRESETDONE,  
    output                              GT_TXPMARESETDONE,
    output                              GT_RXPMARESETDONE,
    output                              GT_TXRESETDONE,
    output                              GT_RXRESETDONE,                 
    
    //--------------------------------------------------------------------------
    //  QPLL Ports
    //--------------------------------------------------------------------------
    input                               GT_QPLL0CLK,
    input                               GT_QPLL0REFCLK,
    input                               GT_QPLL0LOCK,
    input                               GT_QPLL1CLK,
    input                               GT_QPLL1REFCLK,
    input                               GT_QPLL1LOCK,
    
    output      [ 2:0]                  GT_QPLLRATE,
    
    //--------------------------------------------------------------------------
    //  Serial Line Ports
    //--------------------------------------------------------------------------
    input                               GT_RXN,
    input                               GT_RXP,
    
    output                              GT_TXP,
    output                              GT_TXN,
    
    //--------------------------------------------------------------------------
    //  TX Data Ports 
    //--------------------------------------------------------------------------
    input       [63:0]                  GT_TXDATA,
    input       [ 1:0]                  GT_TXDATAK,   
    input                               GT_TXDATA_VALID,
    input                               GT_TXSTART_BLOCK,      
    input       [ 1:0]                  GT_TXSYNC_HEADER,  
    
    //--------------------------------------------------------------------------
    //  RX Data Ports 
    //--------------------------------------------------------------------------
    output      [63:0]                  GT_RXDATA,
    output      [ 1:0]                  GT_RXDATAK,
    output                              GT_RXDATA_VALID,
    output      [ 1:0]                  GT_RXSTART_BLOCK,      
    output      [ 1:0]                  GT_RXSYNC_HEADER,     
    
    //--------------------------------------------------------------------------
    //  PHY Command Ports
    //--------------------------------------------------------------------------
    input                               GT_TXDETECTRX,
    input                               GT_TXELECIDLE,
    input                               GT_TXCOMPLIANCE,
    input                               GT_RXPOLARITY,
    input       [ 1:0]                  GT_POWERDOWN,
    input       [ 1:0]                  GT_RATE,
    input                               GT_RXCDRHOLD,
      
    //--------------------------------------------------------------------------
    //  PHY Status Ports
    //--------------------------------------------------------------------------
    output                              GT_RXVALID,
    output                              GT_PHYSTATUS,
    output                              GT_RXELECIDLE,
    output      [ 2:0]                  GT_RXSTATUS,
      
    //--------------------------------------------------------------------------
    //  TX Equalization Ports 
    //--------------------------------------------------------------------------
    input       [ 2:0]                  GT_TXMARGIN,
    input                               GT_TXSWING,
    input       [ 1:0]                  GT_TXDEEMPH,
    
    //--------------------------------------------------------------------------
    //  TX Equalization Ports (Gen3)
    //--------------------------------------------------------------------------
    input       [ 4:0]                  GT_TXPRECURSOR,
    input       [ 6:0]                  GT_TXMAINCURSOR,
    input       [ 4:0]                  GT_TXPOSTCURSOR,      
    
    //--------------------------------------------------------------------------
    //  PCIe Ports
    //--------------------------------------------------------------------------
    input                               GT_PCIERSTIDLE,        
    input                               GT_PCIERSTTXSYNCSTART, 
    input                               GT_PCIEEQRXEQADAPTDONE,
    input                               GT_PCIEUSERRATEDONE,
             
    output                              GT_PCIEUSERPHYSTATUSRST,    
    output      [ 1:0]                  GT_PCIERATEQPLLPD,                  
    output      [ 1:0]                  GT_PCIERATEQPLLRESET,                
    output                              GT_PCIERATEIDLE,            
    output                              GT_PCIESYNCTXSYNCDONE,                      
    output                              GT_PCIERATEGEN3,    
    output                              GT_PCIEUSERGEN3RDY, 
    output                              GT_PCIEUSERRATESTART,  
                
    //--------------------------------------------------------------------------
    //  USB Ports
    //--------------------------------------------------------------------------
    input                               GT_TXONESZEROS,                        
    input                               GT_RXEQTRAINING,                       
    input                               GT_RXTERMINATION,                        
    
    output                              GT_POWERPRESENT,                                 
                                                          
    //--------------------------------------------------------------------------
    //  TX Sync Alignment Ports
    //--------------------------------------------------------------------------                                                      
    input                               GT_TXSYNCALLIN,
    input                               GT_TXSYNCIN,                                        
                
    output                              GT_TXPHALIGNDONE,            
    output                              GT_TXSYNCOUT,
   
    //--------------------------------------------------------------------------
    //  Loopback & PRBS Ports
    //--------------------------------------------------------------------------     
    input       [ 2:0]                  GT_LOOPBACK,                                              
    input       [ 3:0]                  GT_PRBSSEL,
    input                               GT_TXPRBSFORCEERR, 
    input                               GT_RXPRBSCNTRESET,                                                                                                      

    output                              GT_RXPRBSERR,                                              
    output                              GT_RXPRBSLOCKED,  
      
    //--------------------------------------------------------------------------
    //  GT Status Ports
    //--------------------------------------------------------------------------   
    input                               GT_MASTER_CPLLLOCK,
                                                                                                                      
    output                              GT_CPLLLOCK,
    output                              GT_RXCDRLOCK,
    output                              GT_GEN34_EIOS_DET,
    output                              GT_RXRATEDONE,

    //--------------------------------------------------------------------------
    //  DRP Ports
    //--------------------------------------------------------------------------
    input                               GT_DRPCLK,
    input      [9:0]                    GT_DRPADDR,
    input                               GT_DRPEN,
    input                               GT_DRPWE,
    input      [15:0]                   GT_DRPDI,
    
    output                              GT_DRPRDY,
    output     [15:0]                   GT_DRPDO    
);

//-------------------------------------------------------------------------------------------------
//  Internal Signals
//-------------------------------------------------------------------------------------------------- 
    wire        [127:0]                 txdata;
    wire        [ 15:0]                 txctrl0;
    wire        [ 15:0]                 txctrl1;
    wire        [  7:0]                 txctrl2;
    
    wire        [127:0]                 rxdata;
    wire        [ 15:0]                 rxctrl0;
    
    wire                                pcierategen3;
    wire        [ 15:0]                 pcsrsvdout;
    
    wire                                rxelecidle_int;
    wire                                phy_rxcdrreset;
    wire                                rxcdrreset_int;
 
 
 
    //----------------------------------------------------------------------------------------------
    //  Single vs. Mulit-lane Selection
    //----------------------------------------------------------------------------------------------
    localparam [ 0:0] MULTI_LANE     = (PHY_LANE    == 1) ? 1'b0 : 1'b1;
    localparam [ 0:0] MASTER_LANE    = (GT_LANE_NUM == 0) ? 1'b1 : 1'b0;
    localparam [ 0:0] LOCAL_MASTER   = 1'b1;                                                        // Default for GTH                                      



    //----------------------------------------------------------------------------------------------
    //  PHY Mode
    //----------------------------------------------------------------------------------------------
    localparam        PCS_PCIE_EN = (PHY_MODE == 1) ? "FALSE" : "TRUE";
    localparam [ 0:0] USB_MODE    = (PHY_MODE == 1) ? 1'b1    : 1'b0;



    //----------------------------------------------------------------------------------------------
    //  CPLL_FBDIV - CPLL Feedback (N1) Divider
    //----------------------------------------------------------------------------------------------
    localparam CPLL_FBDIV_45 = (PHY_MAX_SPEED < 3) ? 5 : 4;
    
    
    
    //----------------------------------------------------------------------------------------------
    //  CPLL_FBDIV - CPLL Feedback (N2) Divider
    //----------------------------------------------------------------------------------------------
    localparam CPLL_FBDIV = (PHY_REFCLK_FREQ == 2) ?  2 : 
                            (PHY_REFCLK_FREQ == 1) ?  4 : 5;            
    
    
    
    //----------------------------------------------------------------------------------------------
    // [TX/RX]OUT_DIV - Output Clock Divider
    //----------------------------------------------------------------------------------------------
    localparam OUT_DIV = (PHY_MODE      == 1) ? 1 :
                         (PHY_MAX_SPEED  < 3) ? 2 : 4;  
    
    
    
    //----------------------------------------------------------------------------------------------
    //  [TX/RX]_CLK25_DIV - Clock (25 MHz) Divider
    //----------------------------------------------------------------------------------------------
    localparam CLK25_DIV = (PHY_REFCLK_FREQ == 2) ? 10 : 
                           (PHY_REFCLK_FREQ == 1) ?  5 : 4;
                   
                   
                       
    //----------------------------------------------------------------------------------------------
    //  [TX/RX]_PROGDIV_CFG - Programmable Divider Configuration
    //
    //    Gen1/Gen2 : 250 MHz
    //    Gen3      : 250 or 500 MHz
    //    Gen4      : 500 MHz
    //----------------------------------------------------------------------------------------------
    localparam PROGDIV_CFG = (PHY_MAX_SPEED     < 3) ? 10.0 :                                          
                             (PHY_MAX_SPEED    == 4) ?  4.0 :                                       
                             (PHY_CORECLK_FREQ == 1) ?  8.0 : 4.0;                                 
                       
                       
    
    //----------------------------------------------------------------------------------------------
    //  [TX/RX]PLLCLKSEL - PLL Clock Select   
    //                                                    
    //    2'b00 = CPLL                                                                          
    //    2'b01 = Reserved                                                                          
    //    2'b11 = QPLL0                                                                         
    //    2'b10 = QPLL1                                                                           
    //----------------------------------------------------------------------------------------------
    localparam [ 1:0] PLLCLKSEL = (PHY_MAX_SPEED  < 3) ? 2'b00 : 
                                  (PHY_MAX_SPEED == 3) ? 2'b10 : 2'b11;                                                             
              
                                    
              
    //----------------------------------------------------------------------------------------------
    //  [TX/RX]SYSCLKSEL - System Clock Select   
    //                                                    
    //    2'b00 = CPLL                                                                          
    //    2'b01 = Reserved                                                                          
    //    2'b10 = QPLL0                                                                         
    //    2'b11 = QPLL1                                                                           
    //----------------------------------------------------------------------------------------------                 
    localparam [ 1:0] SYSCLKSEL = (PHY_MAX_SPEED  < 3) ? 2'b00 : 
                                  (PHY_MAX_SPEED == 3) ? 2'b11 : 2'b10;                          
                                  
                                           
                          
     //----------------------------------------------------------------------------------------------
    //  OOBDIVCTL - OOB Divider Control   
    //                                                    
    //    2'd0 = div1                                                                        
    //    2'd1 = div2                                                                        
    //    2'd2 = div4                                                                        
    //    2'd3 = div8                                                                         
    //----------------------------------------------------------------------------------------------                 
    localparam [ 1:0] OOBDIVCTL = (PHY_REFCLK_FREQ == 2) ? 2'd2 : 2'd1; 
                                          
                          
                                                                                                    
    //----------------------------------------------------------------------------------------------
    //  PCIE_PLL_SEL_MODE_GENx - PLL Select Mode for PCIe
    //
    //    2'b00 = CPLL
    //    2'b10 = QPLL0
    //    2'b11 = QPLL1
    //----------------------------------------------------------------------------------------------
    localparam [ 1:0] PCIE_PLL_SEL_MODE_GEN12 = (PHY_MAX_SPEED  < 3) ? 2'b00 : 
                                                (PHY_MAX_SPEED == 3) ? 2'b11 : 2'b10;                 
   
    localparam [ 1:0] PCIE_PLL_SEL_MODE_GEN3  = (PHY_MAX_SPEED  < 3) ? 2'b00 :
                                                (PHY_MAX_SPEED == 3) ? 2'b11 : 2'b10;  
      
    localparam [ 1:0] PCIE_PLL_SEL_MODE_GEN4  = (PHY_MAX_SPEED  < 3) ? 2'b00 :         
                                                (PHY_MAX_SPEED == 3) ? 2'b11 : 2'b10;  
                            
                            
                            
    //----------------------------------------------------------------------------------------------
    //  PCIE_[TX/RX]PMA_CFG - PCIe PMA Configuration    
    //                                         
    //    [   15] : Reserved                                                        
    //    [14:13] : [TX/RX]_INT_DATAWIDTH_G4                                                                    
    //    [12: 9] : [TX/RX]_DATA_WIDTH_G4                                                     
    //    [ 8: 6] : [TX/RX]OUTCLK_DIV_G2                                                        
    //    [ 5: 3] : [TX/RX]OUTCLK_DIV_G3                                                        
    //    [ 2: 0] : [TX/RX]OUTCLK_DIV_G4                                                          
    //----------------------------------------------------------------------------------------------                                                      
    localparam [ 1:0] INT_DATAWIDTH_G4 = 2'd1;
    localparam [ 3:0] DATA_WIDTH_G4    = 4'd4;
    localparam [ 2:0] OUT_DIV_G2       = (PHY_MAX_SPEED  < 3) ? 3'd0 : 3'd1;                                                                                                                                                     
    localparam [ 2:0] OUT_DIV_G3       = (PHY_MAX_SPEED == 4) ? 3'd1 : 3'd0;                                                                                                                                                                    
    localparam [ 2:0] OUT_DIV_G4       = 3'd0;                                                              

    localparam [15:0] PCIE_PMA_CFG = {1'd0,      
                                     INT_DATAWIDTH_G4,                                    
                                     DATA_WIDTH_G4,                                                             
                                     OUT_DIV_G2,                                                 
                                     OUT_DIV_G3,                                                                                              
                                     OUT_DIV_G4};         
    
    
    
    //----------------------------------------------------------------------------------------------
    //  PCIE_BUFG_DIV_CTRL - PCIe BUFG_GT Divider Control
    //
    //    [   15] : BUFG_GT_FSM_CLK
    //    [14:12] : PCLK_DIV_G1
    //    [11:10] : PCLK_DIV_G2  
    //    [ 9: 8] : PCLK_DIV_G3 
    //    [ 7: 6] : PCLK_DIV_G4
    //    [ 5: 0] : Reserved
    //----------------------------------------------------------------------------------------------  
    localparam [ 0:0] BUFG_GT_FSM_CLK    = 1'd0;                                                    // 1'b0 = REFCLK : 1'b1 = PROGDIVCLK
                                                              
    localparam [ 2:0] PCLK_DIV_G1        = (PHY_MODE         == 1) ? 3'd0 :                         // 250 MHz (USB3)
                                           (PHY_MAX_SPEED     < 3) ? 3'd1 :  
                                           (PHY_MAX_SPEED    == 4) ? 3'd3 :                              
                                           (PHY_CORECLK_FREQ == 1) ? 3'd1 : 3'd3;                   // 125 MHz (PCIe)
    
    localparam [ 1:0] PCLK_DIV_G2        = (PHY_MAX_SPEED     < 3) ? 2'd0 : 
                                           (PHY_MAX_SPEED    == 4) ? 2'd1 : 
                                           (PHY_CORECLK_FREQ == 1) ? 2'd0 : 2'd1;                   // 250 MHz
    
    localparam [ 1:0] PCLK_DIV_G3        = PCLK_DIV_G2;                                             // 250 MHz
    
    localparam [ 1:0] PCLK_DIV_G4        = 2'd0;                                                    // 500 MHz
            
    localparam [15:0] PCIE_BUFG_DIV_CTRL = {BUFG_GT_FSM_CLK,                    
                                            PCLK_DIV_G1, 
                                            PCLK_DIV_G2,  
                                            PCLK_DIV_G3,                                                            
                                            PCLK_DIV_G4,
                                            6'd0};
                    
                    
                    
    //----------------------------------------------------------------------------------------------
    //  PCIE_TXPCS_CFG_GEN3 - PCIe TX PCS Configuration
    //                                             
    //    [15:14] : Reserved                                                        
    //    [13:12] : TX_DRIVE_MODE_G3                                                                    
    //    [   11] : ASYNC_EN   
    //    [   10] : TX_XCLK_SEL_G3                                                   
    //    [    9] : TXBUF_EN_G3                                                          
    //    [ 8: 7] : TX_INT_DATAWIDTH_G3
    //    [ 6: 3] : TX_DATA_WIDTH_G3
    //    [    2] : TX_SYNC_MODE
    //    [    1] : DRP_EXT_CTRL                                                         
    //    [    0] : Reserved                                                         
    //----------------------------------------------------------------------------------------------                                                      
    localparam [ 1:0] TX_DRIVE_MODE_G3    = 2'd2;                                      // "PIPEGEN3"
    localparam [ 0:0] ASYNC_EN            = (PHY_REFCLK_MODE != 0) ? 1'd1 : 1'd0;      // 1'b0 = Async : 1'b1 = Sync
    localparam [ 0:0] TX_XCLK_SEL_G3      = 1'd1;                                      // "TXUSER" when bypassing TX buffer                                                                                                                                                     
    localparam [ 0:0] TXBUF_EN_G3         = 1'd0;                                      // "FALSE"                                                                                                                                        
    localparam [ 1:0] TX_INT_DATAWIDTH_G3 = 2'd1;                                      //  4-byte
    localparam [ 3:0] TX_DATA_WIDTH_G3    = 4'd4;                                      // 32-bit 
    localparam [ 0:0] TX_SYNC_MODE        = 1'd1;                                      // Auto 
    localparam [ 0:0] DRP_EXT_CTRL        = 1'd0;                                      // Disable (Advance feature) 
    
    localparam [15:0] PCIE_TXPCS_CFG_GEN3 = {2'd0,
                                             TX_DRIVE_MODE_G3,
                                             ASYNC_EN,
                                             TX_XCLK_SEL_G3,
                                             TXBUF_EN_G3,
                                             TX_INT_DATAWIDTH_G3,
                                             TX_DATA_WIDTH_G3,
                                             TX_SYNC_MODE,
                                             DRP_EXT_CTRL,
                                             1'd0};
    
    
    
    //----------------------------------------------------------------------------------------------
    //  PCIE_RXPCS_CFG_GEN3 - PCIe RX PCS Configuration  
    //                                                                                                  
    //    [   15] : RX_DFE_LPM_HOLD_DURING_EIDLE_G3                                                                 
    //    [   14] : RXCDR_PH_RESET_ON_EIDLE_G3  
    //    [   13] : RXCDR_FR_RESET_ON_EIDLE_G3                                             
    //    [   12] : RXCDR_HOLD_DURING_EIDLE_G3                                                      
    //    [   11] : CLK_CORRECT_USE_G3
    //    [   10] : RX_XCLK_SEL_G3
    //    [    9] : RXBUF_EN_G3
    //    [ 8: 7] : RX_INT_DATA_WIDTH_G3
    //    [ 6: 3] : RX_DATA_WIDTH_G3
    //    [    2] : RX_SYNC_MODE                                                        
    //    [    1] : RATE_FSM_CLK  
    //    [    0] : RXVALID_GATE_G3                                                
    //----------------------------------------------------------------------------------------------                                                      
    localparam [ 0:0] RX_DFE_LPM_HOLD_DURING_EIDLE_G3 = 1'd0;                          // 
    localparam [ 0:0] RXCDR_PH_RESET_ON_EIDLE_G3      = 1'd0;                          // 
    localparam [ 0:0] RXCDR_FR_RESET_ON_EIDLE_G3      = 1'd0;                          //                                                                                                                                          
    localparam [ 0:0] RXCDR_HOLD_DURING_EIDLE_G3      = 1'd0;                          //             
    localparam [ 0:0] CLK_CORRECT_USE_G3              = 1'd1;                          // "TRUE"       
    localparam [ 0:0] RX_XCLK_SEL_G3                  = 1'd0;                          // "RXDES" when using RX buffer                                                                              
    localparam [ 0:0] RXBUF_EN_G3                     = 1'd1;                          // "TRUE"
    localparam [ 1:0] RX_INT_DATA_WIDTH_G3            = 2'd1;                          //  4-byte  
    localparam [ 3:0] RX_DATA_WIDTH_G3                = 4'd4;                          // 32-bit  
    localparam [ 0:0] RX_SYNC_MODE                    = 1'd1;                          // Auto
    localparam [ 0:0] RATE_FSM_CLK                    = 1'd0;                          // 1'b0 = REFCLK : 1'b1 = PCLK
    localparam [ 0:0] RXVALID_GATE_G3                 = 1'd1;
    
    localparam [15:0] PCIE_RXPCS_CFG_GEN3 = {RX_DFE_LPM_HOLD_DURING_EIDLE_G3,
                                             RXCDR_PH_RESET_ON_EIDLE_G3,
                                             RXCDR_FR_RESET_ON_EIDLE_G3,
                                             RXCDR_HOLD_DURING_EIDLE_G3,
                                             CLK_CORRECT_USE_G3,
                                             RX_XCLK_SEL_G3,
                                             RXBUF_EN_G3,
                                             RX_INT_DATA_WIDTH_G3,
                                             RX_DATA_WIDTH_G3,
                                             RX_SYNC_MODE,
                                             RATE_FSM_CLK,
                                             RXVALID_GATE_G3};
    
    //----------------------------------------------------------------------------------------------
    //  PCIe CDR for Gen1/Gen2
    //  USB CDR for Gen1 (5G) uses same setting
    //----------------------------------------------------------------------------------------------   
    localparam [15:0] RXCDR_CFG0      = 16'b0000_0000_0000_0010;
    localparam [15:0] RXCDR_CFG1      = 16'b0000_0000_0000_0000;
    localparam [15:0] RXCDR_CFG2      = (PHY_REFCLK_MODE == 2) ? 16'b0000_0001_1110_0100 : 16'b0000001001011001;
    localparam [15:0] RXCDR_CFG3      = 16'b0000_0000_0001_0010; 
    localparam [15:0] RXCDR_CFG4      = 16'b0101_1100_1111_0110;
    localparam [15:0] RXCDR_CFG5      = 16'b1011_0100_0110_1011;
    
    //----------------------------------------------------------------------------------------------
    //  PCIe CDR for Gen3
    //---------------------------------------------------------------------------------------------- 
    localparam [15:0] RXCDR_CFG0_GEN3 = RXCDR_CFG0;
    localparam [15:0] RXCDR_CFG1_GEN3 = RXCDR_CFG1;
    localparam [15:0] RXCDR_CFG2_GEN3 = (PHY_REFCLK_MODE == 2) ? 16'b0000_0000_0011_0110 : 16'b0000_0000_0011_0100;
    localparam [15:0] RXCDR_CFG3_GEN3 = RXCDR_CFG3; 
    localparam [15:0] RXCDR_CFG4_GEN3 = RXCDR_CFG4;
    localparam [15:0] RXCDR_CFG5_GEN3 = 16'b0001_0100_0110_1011;
    
    //----------------------------------------------------------------------------------------------
    //  PCIe CDR for Gen4
    //---------------------------------------------------------------------------------------------- 
    localparam [15:0] RXCDR_CFG2_GEN4 = (PHY_REFCLK_MODE == 2) ? 16'b0000_0000_0100_0110 : 16'b0000_0000_0011_0100;          
    localparam [15:0] RXCDR_CFG3_GEN4 = RXCDR_CFG4_GEN3;

    //----------------------------------------------------------------------------------------------
    //  PCIe RX Buffer for Gen1/Gen2
    //----------------------------------------------------------------------------------------------  
    localparam [5:0] PCIE_CLK_COR_MAX_LAT     = (PHY_REFCLK_MODE == 2) ? 6'd28 : (PHY_REFCLK_MODE == 1) ? 6'd20 : 6'd20;
    localparam [5:0] PCIE_CLK_COR_MIN_LAT     = (PHY_REFCLK_MODE == 2) ? 6'd22 : (PHY_REFCLK_MODE == 1) ? 6'd17 : 6'd4;
    localparam [5:0] PCIE_RXBUF_THRESH_OVFLW  = (PHY_REFCLK_MODE == 2) ? 6'd63 : (PHY_REFCLK_MODE == 1) ? 6'd31 : 6'd31;
    localparam [5:0] PCIE_RXBUF_THRESH_UNDFLW = (PHY_REFCLK_MODE == 2) ? 6'd8  : (PHY_REFCLK_MODE == 1) ? 6'd8  : 6'd1;
    
    //----------------------------------------------------------------------------------------------
    //  PCIe RX Buffer for Gen3/Gen4
    //----------------------------------------------------------------------------------------------  
    localparam [4:0] PCIE3_CLK_COR_EMPTY_THRSH = 5'd0;
    localparam [5:0] PCIE3_CLK_COR_FULL_THRSH  = (PHY_REFCLK_MODE == 2) ? 6'd32 : (PHY_REFCLK_MODE == 1) ? 6'd16 : 6'd16;
    localparam [4:0] PCIE3_CLK_COR_MAX_LAT     = (PHY_REFCLK_MODE == 2) ? 5'd16 : (PHY_REFCLK_MODE == 1) ? 5'd8  : 5'd4;
    localparam [4:0] PCIE3_CLK_COR_MIN_LAT     = (PHY_REFCLK_MODE == 2) ? 5'd12 : (PHY_REFCLK_MODE == 1) ? 5'd4  : 5'd0;
    localparam [5:0] PCIE3_CLK_COR_THRSH_TIMER = (PHY_REFCLK_MODE == 2) ? 6'd4  : (PHY_REFCLK_MODE == 1) ? 6'd8  : 6'd8;
    
    //----------------------------------------------------------------------------------------------
    //  TX Electrical Idle Attributes for USB3 and PCIe
    //---------------------------------------------------------------------------------------------- 
    localparam [ 2:0]  TX_EIDLE_ASSERT_DELAY   = (PHY_MODE == 1)      ? 3'd0 :
                                                 (PHY_MAX_SPEED == 4) ? 3'd6 :   // For PCIe Gen4 EIOS TX
                                                                        3'd5 ;   // For PCIe Gen3 EIOS TX    
    localparam [ 2:0]  TX_EIDLE_DEASSERT_DELAY = (PHY_MODE == 1) ? 3'd1 : 3'd3;
    
    //----------------------------------------------------------------------------------------------
    //  Comma Align and Detect Attributres for USB3 and PCIe                                                                  
    //----------------------------------------------------------------------------------------------     
    localparam         ALIGN_COMMA_DOUBLE  = (PHY_MODE == 1) ? "TRUE" : "FALSE";                      
    localparam         SHOW_REALIGN_COMMA  = (PHY_MODE == 1) ? "TRUE" : "FALSE";  
    
    //----------------------------------------------------------------------------------------------
    //  Clock Correction Attributes for USB3 and PCIe
    //----------------------------------------------------------------------------------------------
    localparam [ 5:0]  CLK_COR_MAX_LAT      = (PHY_MODE == 1) ?  6'd16        : PCIE_CLK_COR_MAX_LAT;
    localparam [ 5:0]  CLK_COR_MIN_LAT      = (PHY_MODE == 1) ?  6'd13        : PCIE_CLK_COR_MIN_LAT;
    localparam         CLK_COR_KEEP_IDLE    = (PHY_MODE == 1) ? "FALSE"       : "TRUE";
    localparam [ 9:0]  CLK_COR_SEQ_1_1      = (PHY_MODE == 1) ? 10'b100111100 : 10'b0100011100;
    localparam [ 9:0]  CLK_COR_SEQ_1_2      = (PHY_MODE == 1) ? 10'b100111100 : 10'b0000000000;
    localparam [ 3:0]  CLK_COR_SEQ_2_ENABLE = (PHY_MODE == 1) ?  4'b0000      :  4'b1111;
    localparam [ 1:0]  CLK_COR_SEQ_LEN      = (PHY_MODE == 1) ? 2             : 1;

    //----------------------------------------------------------------------------------------------
    //  RX Buffer Attributes for USB3 and PCIe                                                                  
    //----------------------------------------------------------------------------------------------
    localparam [ 5:0]  RXBUF_THRESH_OVFLW  = (PHY_MODE == 1) ? 32 : PCIE_RXBUF_THRESH_OVFLW;                                                            
    localparam [ 5:0]  RXBUF_THRESH_UNDFLW = (PHY_MODE == 1) ?  6 : PCIE_RXBUF_THRESH_UNDFLW;                                    
    
    //----------------------------------------------------------------------------------------------
    //  RX Common Mode Select for USB3 and PCIe        
    //
    //    0 = AVTT
    //    1 = GND
    //    2 = Floating
    //    3 = Programmable                                                         
    //----------------------------------------------------------------------------------------------
    localparam integer RX_CM_SEL = (PHY_MODE == 1) ?  1 : 3;   
   
    //----------------------------------------------------------------------------------------------
    //  GT Attributes for USB3 and PCIe                                                                  
    //----------------------------------------------------------------------------------------------  
    localparam         SIM_TX_EIDLE_DRIVE_LEVEL = (PHY_MODE == 1) ? "Z"   : "LOW";    
    localparam         RXSLIDE_MODE             = (PHY_MODE == 1) ? "OFF" : "PMA";   

    //----------------------------------------------------------------------------------------------
    //  Reserved Attributes for USB3 and PCIe                                                                  
    //----------------------------------------------------------------------------------------------      
    localparam [ 8:0]  USB_LFPS_DET      = (PHY_REFCLK_FREQ == 0) ? 9'b011001001 : 9'b011001010; 
    localparam         RXTERMINATION_DRP = 1'd1;
    localparam [ 1:0]  RX_CM_SEL_USB     = 2'd3;
    
    localparam [15:0]  PCS_RSVD0         = {USB_LFPS_DET, 4'd0, RXTERMINATION_DRP, RX_CM_SEL_USB};
        
    //----------------------------------------------------------------------------------------------
    //  Other Attributes based on latest 2015.3 rules                                                                 
    //----------------------------------------------------------------------------------------------   
    localparam [3:0]   RX_SUM_VCMTUNE    = (PHY_MODE         == 1) ? 4'b0110 : 
                                           (PHY_MAX_SPEED     < 3) ? 4'b0110 : 4'b1010; 
                                           
    localparam [3:0]   RX_SUM_IREF_TUNE  = (PHY_MODE         == 1) ? 4'b0100 : 
                                           (PHY_MAX_SPEED     < 3) ? 4'b0100 : 4'b1001; 
                                           
    localparam         RXDFE_PWR_SAVING  = (PHY_MODE         == 1) ? 1'b0 :
                                           (PHY_MAX_SPEED    == 4) ? 1'b1 : 1'b0;
                                           
    localparam         TX_PI_BIASSET     = (PHY_MODE         == 1) ? 0 :
                                           (PHY_MAX_SPEED     < 3) ? 0 :
                                           (PHY_MAX_SPEED    == 3) ? 1 : 3;
    
    localparam  [15:0] RXPI_CFG0         = (PHY_MODE         == 1) ? 16'h1200 :
                                           (PHY_MAX_SPEED     < 3) ? 16'h1200 :
                                           (PHY_MAX_SPEED    == 3) ? 16'h2202 : 16'b0000000100000100;
//--------------------------------------------------------------------------------------------------
//  GT Channel
//--------------------------------------------------------------------------------------------------
generate
  if (PHY_GT_XCVR == "GTY" || PHY_GT_XCVR == "GTY64") begin: GTY_CHANNEL
//--------------------------------------------------------------------------------------------------
//  GTY Channel
//--------------------------------------------------------------------------------------------------
GTYE4_CHANNEL #
(  
    //----------------------------------------------------------------------------------------------
    //  Simulation Attributes
    //----------------------------------------------------------------------------------------------
    .SIM_MODE                           ("FAST"),                                    
    .SIM_RECEIVER_DETECT_PASS           ("TRUE"),
    .SIM_RESET_SPEEDUP                  ("TRUE"),
    .SIM_TX_EIDLE_DRIVE_LEVEL           (SIM_TX_EIDLE_DRIVE_LEVEL),
    //.SIM_VERSION                        (1),                             
   
    //----------------------------------------------------------------------------------------------     
    //  Clock Attributes
    //----------------------------------------------------------------------------------------------                       
    .TXREFCLKDIV2_SEL                   ( 1'b0),                              
    .RXREFCLKDIV2_SEL                   ( 1'b0),                                
    .TX_CLK25_DIV                       (CLK25_DIV),                                                    
    .RX_CLK25_DIV                       (CLK25_DIV),                                                    
    .TX_CLKMUX_EN                       ( 1'b1),                                                
    .RX_CLKMUX_EN                       ( 1'b1),                                                
    .TX_XCLK_SEL                        ("TXUSR"),                                              
    .RX_XCLK_SEL                        ("RXDES"),   
    .TXOUT_DIV                          (OUT_DIV), 
    .RXOUT_DIV                          (OUT_DIV), 
    .LOCAL_MASTER                       (LOCAL_MASTER),   
    .RX_CLK_SLIP_OVRD                   ( 5'b00000),  
    .RXPMACLK_SEL                       ("DATA"),                                                                                                                           
    .USE_PCS_CLK_PHASE_SEL              ( 1'b0),           
   
    //----------------------------------------------------------------------------------------------     
    //  Programmable Divider Attributes
    //----------------------------------------------------------------------------------------------                                                                                                                       
    .TX_PROGCLK_SEL                     ("CPLL"),                               
    .TX_PROGDIV_CFG                     (PROGDIV_CFG),                      
    .RX_PROGDIV_CFG                     (PROGDIV_CFG),   
    .TX_PROGDIV_RATE                    (16'h0001),                          
    .RX_PROGDIV_RATE                    (16'h0001),                                   
               
    //----------------------------------------------------------------------------------------------
    //  CPLL Attributes
    //----------------------------------------------------------------------------------------------                 
    .CPLL_CFG0                          (16'h0000), //(16'h20FA),                             // Optimize for PCIe PLL compliance   [Changed for extracted model]
    .CPLL_CFG1                          (16'h81E4), //(16'h24AA),               [Changed for extracted model]
    .CPLL_CFG2                          (16'hF007),                             
    .CPLL_CFG3                          ( 6'h00),  
    .CPLL_FBDIV                         (CPLL_FBDIV),  
    .CPLL_FBDIV_45                      (CPLL_FBDIV_45),    
    .CPLL_INIT_CFG0                     (16'h001E),                
    .CPLL_LOCK_CFG                      (16'h01EC), //(16'h01E8),                             // Bit[0] must be LOW   [Changed for extracted model]
    .CPLL_REFCLK_DIV                    ( 1),     
             
    //----------------------------------------------------------------------------------------------
    //  Reset Attributes
    //----------------------------------------------------------------------------------------------                
    //.RESET_POWERSAVE_DISABLE            ( 1'b0),   
                                                                              
    //----------------------------------------------------------------------------------------------
    //  Reset Time Attributes
    //----------------------------------------------------------------------------------------------    
    .TX_DIVRESET_TIME                   ( 5'b00001),
    .TXPCSRESET_TIME	                ( 5'b00001),
    .TXPMARESET_TIME	                ( 5'b00001),
    .RX_DIVRESET_TIME                   ( 5'b00001),
    .RXBUFRESET_TIME                    ( 5'b00001),
    .RXCDRFREQRESET_TIME                ( 5'b10000), //( 5'b00001),  [Changed for extracted model]
    .RXCDRPHRESET_TIME                  ( 5'b00001),    
    .RXDFELPMRESET_TIME                 ( 7'b0001111),    
    .RXISCANRESET_TIME	                ( 5'b00001), 
    .RXOSCALRESET_TIME	                ( 5'b00011), 
    .RXPCSRESET_TIME	                  ( 5'b00001),   
    .RXPMARESET_TIME	                  ( 5'b00001),   
               
    //----------------------------------------------------------------------------------------------
    //  PCIe Attributes
    //----------------------------------------------------------------------------------------------
    .PCIE_GEN4_64BIT_INT_EN             (PHY_GEN4_64BIT_EN),  // THIS ATTRIBUTE IS NEW AND MAY NOT BE AVAILABLE IN EARLY GT MODELS
    .PCIE_BUFG_DIV_CTRL                 (PCIE_BUFG_DIV_CTRL),                  
    .PCIE_RXPCS_CFG_GEN3                (PCIE_RXPCS_CFG_GEN3),                 
    .PCIE_RXPMA_CFG                     (PCIE_PMA_CFG),                        
    .PCIE_TXPCS_CFG_GEN3                (PCIE_TXPCS_CFG_GEN3),                 
    .PCIE_TXPMA_CFG                     (PCIE_PMA_CFG),                        
    .PCS_PCIE_EN                        (PCS_PCIE_EN),  
    .PCIE_PLL_SEL_MODE_GEN12            (PCIE_PLL_SEL_MODE_GEN12),                  
    .PCIE_PLL_SEL_MODE_GEN3             (PCIE_PLL_SEL_MODE_GEN3),  
    .PCIE_PLL_SEL_MODE_GEN4             (PCIE_PLL_SEL_MODE_GEN4),

    //---------------------------------------------------------------------------------------------- 
    //  Data Width Attributes
    //----------------------------------------------------------------------------------------------                          
    .TX_DATA_WIDTH                      (20),                                                                                                                                         
    .RX_DATA_WIDTH                      (20),  
    .TX_INT_DATAWIDTH                   ( 0),                                                                
    .RX_INT_DATAWIDTH                   ( 0),   
    .TX_FABINT_USRCLK_FLOP              ( 1'b0), 
    .RX_FABINT_USRCLK_FLOP              ( 1'b0),                                                    
              
    //----------------------------------------------------------------------------------------------
    //  Analog Front End Attributes
    //----------------------------------------------------------------------------------------------
    .LPBK_BIAS_CTRL	                    ( 3'b000),                           
    .LPBK_EN_RCAL_B	                    ( 1'b0),                             
    .LPBK_EXT_RCAL	                    ( 4'b0000),                          
    .LPBK_RG_CTRL	                      ( 4'b0000),                             
    .RX_AFE_CM_EN                       ( 1'b0),
    .RX_BIAS_CFG0                       (16'h1534),
    .RX_CM_BUF_CFG                      ( 4'b1010),
    .RX_CM_BUF_PD                       ( 1'b0),                                           
    .RX_CM_SEL                          (RX_CM_SEL),                                                        
    .RX_CM_TRIM                         (10),    
    .RX_TUNE_AFE_OS                     ( 2'b00),
    .TERM_RCAL_CFG                      (15'b100001000010000),                                     
    .TERM_RCAL_OVRD                     ( 3'b000),             
                                                                                                    
    //----------------------------------------------------------------------------------------------  
    //  Receiver Detection Attributes
    //----------------------------------------------------------------------------------------------                                      
    .TX_RXDETECT_CFG                    (14'h0032),                                                      
    .TX_RXDETECT_REF                    (3),                                  
    
    //----------------------------------------------------------------------------------------------  
    //  TX Electrical Idle Attributes
    //----------------------------------------------------------------------------------------------   
    .TX_EIDLE_ASSERT_DELAY              (TX_EIDLE_ASSERT_DELAY),                            
    .TX_EIDLE_DEASSERT_DELAY            (TX_EIDLE_DEASSERT_DELAY),             
    .TX_IDLE_DATA_ZERO                  ( 1'b0),                                // Optimized for PCIe      
 
    //----------------------------------------------------------------------------------------------  
    //  RX OOB Attributes
    //----------------------------------------------------------------------------------------------   
    .OOB_PWRUP                          ( 1'b1),                                
    .OOBDIVCTL                          (OOBDIVCTL),                                            
    .RX_SIG_VALID_DLY                   ( 4),                                   // Optimized for PCIe
    .RXOOB_CFG                          ( 9'b000000110),                          
    .RXOOB_CLK_CFG                      ("PMA"),      
    
    //----------------------------------------------------------------------------------------------  
    //  RX Electrical Idle Attributes
    //----------------------------------------------------------------------------------------------                                                   
    .RX_DFE_LPM_HOLD_DURING_EIDLE       ( 1'b0),                                
    .RXBUF_EIDLE_HI_CNT                 ( 4'b0100),                             // Optimized for PCIe
    .RXBUF_EIDLE_LO_CNT                 ( 4'b0000),
    .RXBUF_RESET_ON_EIDLE               ("TRUE"),
    .RXCDR_FR_RESET_ON_EIDLE            ( 1'b0),
    .RXCDR_PH_RESET_ON_EIDLE            ( 1'b0),
    .RXCDR_HOLD_DURING_EIDLE            ( 1'b0),                                // Optimized for PCIe
    .RXELECIDLE_CFG                     ("SIGCFG_1"),                           // Optimized for PCIe
 
    //----------------------------------------------------------------------------------------------  
    //  Power Down Attributes
    //----------------------------------------------------------------------------------------------   
    .PD_TRANS_TIME_FROM_P2              (12'h03C),                                                     
    .PD_TRANS_TIME_NONE_P2              ( 8'h19),                                                      
    .PD_TRANS_TIME_TO_P2                ( 8'h64),   
    .TX_PMA_POWER_SAVE                  ( 1'b0),   
    .RX_PMA_POWER_SAVE                  ( 1'b0),                               
  
    //----------------------------------------------------------------------------------------------  
    //  Rate Change Attributes
    //---------------------------------------------------------------------------------------------- 
    .RATE_SW_USE_DRP                    ( 1'b0),                                // Advance PCIe feature
    .TRANS_TIME_RATE                    ( 8'h0E),             
    .TXBUF_RESET_ON_RATE_CHANGE         ("TRUE"),                              
    .RXBUF_RESET_ON_RATE_CHANGE         ("TRUE"),                              

    //----------------------------------------------------------------------------------------------
    //  TX Driver Attributes
    //----------------------------------------------------------------------------------------------                                   
    .TX_DEEMPH0                         ( 6'b010100),                           // -6.0 dB 
    .TX_DEEMPH1                         ( 6'b001101),                           // -3.5 dB
    .TX_DEEMPH2                         ( 6'b000000),                           //  0.0 dB 
    .TX_DEEMPH3                         ( 6'b000000),                           //  0.0 dB  
    .TX_DRIVE_MODE                      ("PIPE"),                                
    .TX_LOOPBACK_DRIVE_HIZ              ("FALSE"),                   
    .TX_MAINCURSOR_SEL                  ( 1'b0),   
    .TX_MARGIN_FULL_0                   ( 7'b1001111),                          // 1200 mV
    .TX_MARGIN_FULL_1                   ( 7'b1001110),                          // 1100 mV
    .TX_MARGIN_FULL_2                   ( 7'b1001100),                          // 1000 mV 
    .TX_MARGIN_FULL_3                   ( 7'b1001010),                          //  900 mV
    .TX_MARGIN_FULL_4                   ( 7'b1001000),                          //  800 mV
    .TX_MARGIN_LOW_0                    ( 7'b1000110),                          //  700 mV            
    .TX_MARGIN_LOW_1                    ( 7'b1000101),                          //  600 mV           
    .TX_MARGIN_LOW_2                    ( 7'b1000011),                          //  500 mV          
    .TX_MARGIN_LOW_3                    ( 7'b1000010),                          //  400 mV           
    .TX_MARGIN_LOW_4                    ( 7'b1000000),                          //  300 mV                               
   
    //----------------------------------------------------------------------------------------------    
    //  Comma Align & Detect Attributes
    //----------------------------------------------------------------------------------------------       
    .ALIGN_COMMA_DOUBLE                 (ALIGN_COMMA_DOUBLE),                                                  
    .ALIGN_COMMA_ENABLE                 (10'b1111111111),                                           
    .ALIGN_COMMA_WORD                   ( 1),                                                       
    .ALIGN_MCOMMA_DET                   ("TRUE"),                                                   
    .ALIGN_MCOMMA_VALUE                 (10'b1010000011),                                           
    .ALIGN_PCOMMA_DET                   ("TRUE"),                                                   
    .ALIGN_PCOMMA_VALUE                 (10'b0101111100),                                           
    .DEC_MCOMMA_DETECT                  ("TRUE"),                                                      
    .DEC_PCOMMA_DETECT                  ("TRUE"),                                                      
    .DEC_VALID_COMMA_ONLY               ("FALSE"),                                                     
    .SHOW_REALIGN_COMMA                 (SHOW_REALIGN_COMMA),       
   
    //----------------------------------------------------------------------------------------------   
    //  8B/10B Attributes                                                                             
    //----------------------------------------------------------------------------------------------                   
    .RX_DISPERR_SEQ_MATCH               ("TRUE"),        
   
    //----------------------------------------------------------------------------------------------  
    //  TX Buffer Attributes
    //----------------------------------------------------------------------------------------------                      
    .TX_FIFO_BYP_EN                     ( 1'b1),                                
    .TXBUF_EN                           ("FALSE"),        
    .TXFIFO_ADDR_CFG                    ("LOW"),                                                                                      
 
    //----------------------------------------------------------------------------------------------
    //  RX Buffer Attributes                                                                        
    //----------------------------------------------------------------------------------------------     
    .RXBUF_ADDR_MODE                    ("FULL"),                               
    .RXBUF_EN                           ("TRUE"),
    .RXBUF_RESET_ON_CB_CHANGE           ("TRUE"),
    .RXBUF_RESET_ON_COMMAALIGN          ("FALSE"),
    .RXBUF_THRESH_OVFLW                 (RXBUF_THRESH_OVFLW),                                                      
    .RXBUF_THRESH_OVRD                  ("TRUE"),                             
    .RXBUF_THRESH_UNDFLW                (RXBUF_THRESH_UNDFLW),                                    
    .RX_BUFFER_CFG                      ( 6'b000000),
    .RX_DEFER_RESET_BUF_EN              ("TRUE"), 
   
    //----------------------------------------------------------------------------------------------   
    //  PCIe Gen3 RX Buffer Attributes                                                                                   
    //----------------------------------------------------------------------------------------------   
    .PCI3_AUTO_REALIGN                  ("OVR_1K_BLK"),                           
    .PCI3_PIPE_RX_ELECIDLE              ( 1'b0),                                
    .PCI3_RX_ASYNC_EBUF_BYPASS          ( 2'b00),                               
    .PCI3_RX_ELECIDLE_EI2_ENABLE        ( 1'b0),                                
    .PCI3_RX_ELECIDLE_H2L_COUNT         ( 6'b000000),                           
    .PCI3_RX_ELECIDLE_H2L_DISABLE       ( 3'b000),                              
    .PCI3_RX_ELECIDLE_HI_COUNT          ( 6'b000000),                           
    .PCI3_RX_ELECIDLE_LP4_DISABLE       ( 1'b0),                                
    .PCI3_RX_FIFO_DISABLE               ( 1'b0),                                
       
    //----------------------------------------------------------------------------------------------   
    //  PCIe Gen3 Clock Correction Attributes                                                                                   
    //----------------------------------------------------------------------------------------------          
    .PCIE3_CLK_COR_EMPTY_THRSH             (PCIE3_CLK_COR_EMPTY_THRSH),                           
    .PCIE3_CLK_COR_FULL_THRSH              (PCIE3_CLK_COR_FULL_THRSH),                          
    .PCIE3_CLK_COR_MAX_LAT                 (PCIE3_CLK_COR_MAX_LAT),                          
    .PCIE3_CLK_COR_MIN_LAT                 (PCIE3_CLK_COR_MIN_LAT),                          
    .PCIE3_CLK_COR_THRSH_TIMER             (PCIE3_CLK_COR_THRSH_TIMER),                      
       
    //---------------------------------------------------------------------------------------------- 
    //  Clock Correction Attributes
    //----------------------------------------------------------------------------------------------             
    .CBCC_DATA_SOURCE_SEL               ("DECODED"),  
    .CLK_COR_KEEP_IDLE                  (CLK_COR_KEEP_IDLE),
    .CLK_COR_MAX_LAT                    (CLK_COR_MAX_LAT),                                   
    .CLK_COR_MIN_LAT                    (CLK_COR_MIN_LAT),                                  
    .CLK_COR_PRECEDENCE                 ("TRUE"),
    .CLK_COR_REPEAT_WAIT                (0),
    .CLK_COR_SEQ_1_1                    (CLK_COR_SEQ_1_1),
    .CLK_COR_SEQ_1_2                    (CLK_COR_SEQ_1_2),
    .CLK_COR_SEQ_1_3                    (10'b0000000000),
    .CLK_COR_SEQ_1_4                    (10'b0000000000),
    .CLK_COR_SEQ_1_ENABLE               (4'b1111),
    .CLK_COR_SEQ_2_1                    (10'b0000000000),
    .CLK_COR_SEQ_2_2                    (10'b0000000000),
    .CLK_COR_SEQ_2_3                    (10'b0000000000),
    .CLK_COR_SEQ_2_4                    (10'b0000000000),
    .CLK_COR_SEQ_2_ENABLE               (CLK_COR_SEQ_2_ENABLE),
    .CLK_COR_SEQ_2_USE                  ("FALSE"),
    .CLK_COR_SEQ_LEN                    (CLK_COR_SEQ_LEN),
    .CLK_CORRECT_USE                    ("TRUE"),                
       
    //---------------------------------------------------------------------------------------------- 
    //  FTS Deskew Attributes                                                                            
    //----------------------------------------------------------------------------------------------                                         
    .FTS_DESKEW_SEQ_ENABLE              ( 4'b1111),                                        
    .FTS_LANE_DESKEW_CFG                ( 4'b1111),                                          
    .FTS_LANE_DESKEW_EN                 ("FALSE"),           
       
    //---------------------------------------------------------------------------------------------- 
    //  Channel Bonding Attributes (Disabled)
    //----------------------------------------------------------------------------------------------          
    .CHAN_BOND_KEEP_ALIGN               ("FALSE"),
    .CHAN_BOND_MAX_SKEW                 ( 1),
    .CHAN_BOND_SEQ_1_1                  (10'b0000000000),
    .CHAN_BOND_SEQ_1_2                  (10'b0000000000),
    .CHAN_BOND_SEQ_1_3                  (10'b0000000000),
    .CHAN_BOND_SEQ_1_4                  (10'b0000000000),
    .CHAN_BOND_SEQ_1_ENABLE             ( 4'b1111),
    .CHAN_BOND_SEQ_2_1                  (10'b0000000000),
    .CHAN_BOND_SEQ_2_2                  (10'b0000000000),
    .CHAN_BOND_SEQ_2_3                  (10'b0000000000),
    .CHAN_BOND_SEQ_2_4                  (10'b0000000000),  
    .CHAN_BOND_SEQ_2_ENABLE             ( 4'b1111),
    .CHAN_BOND_SEQ_2_USE                ("FALSE"), 
    .CHAN_BOND_SEQ_LEN                  ( 1),                                                           
  
    //----------------------------------------------------------------------------------------------            
    //  TX Sync Alignment Attributes                                                                              
    //----------------------------------------------------------------------------------------------     
    .TXDLY_CFG                          (16'b0000000000011111),    
    .TXDLY_LCFG                         (16'b0000000001010000),                
    .TXPH_CFG                           (16'b0000000100000011),
    .TXPH_CFG2                          (16'b0000000000000000),                 
    .TXPH_MONITOR_SEL                   ( 5'b00000),
    .TXPHDLY_CFG0                       (16'b0110000000100000),                 
    .TXPHDLY_CFG1                       (16'b0000000000000010),              
                                                                                    
    //----------------------------------------------------------------------------------------------            
    //  TX Auto Sync Alignment Attributes                                                                               
    //----------------------------------------------------------------------------------------------                
    .TXSYNC_MULTILANE                   (MULTI_LANE),                                                                                                              
    .TXSYNC_OVRD                        (1'b0),                                 // Select auto TXSYNC mode                                                                                 
    .TXSYNC_SKIP_DA                     (1'b0),                     
                                                                                                    
    //----------------------------------------------------------------------------------------------            
    //  RX Sync Alignment Attributes (Not used)                                                                             
    //----------------------------------------------------------------------------------------------    
  //.RXDLY_CFG                          (16'h001F),   
  //.RXDLY_LCFG                         (16'h0030),   
  //.RXPH_MONITOR_SEL                   (5'b00000),
  //.RXPHBEACON_CFG                     (16'h0000),
  //.RXPHDLY_CFG                        (16'h2020),
  //.RXPHSAMP_CFG                       (16'h2100),
  //.RXPHSLIP_CFG                       (16'h9933),                             
     
    //----------------------------------------------------------------------------------------------            
    //  RX Auto Sync Alignment Attributes (Not used)                                                                                
    //----------------------------------------------------------------------------------------------                
  //.RXSYNC_MULTILANE                   (1'b0),                                                                                                              
  //.RXSYNC_OVRD                        (1'b0),                                                                                         
  //.RXSYNC_SKIP_DA                     (1'b0),                   
  
    //----------------------------------------------------------------------------------------------  
    //  Gearbox Attributes (Not used)                                                                
    //---------------------------------------------------------------------------------------------- 
  //.GEARBOX_MODE                       ( 5'b00000), 
  //.TX_SAMPLE_PERIOD                   ( 3'b101),
  //.RX_SAMPLE_PERIOD                   ( 3'b101),
  //.TXGEARBOX_EN                       ("FALSE"),
  //.RXGEARBOX_EN                       ("FALSE"),    
  //.TXGBOX_FIFO_INIT_RD_ADDR           ( 4),
  //.RXGBOX_FIFO_INIT_RD_ADDR           ( 4),
  //.RXSLIDE_AUTO_WAIT                  ( 7),                                                         
    .RXSLIDE_MODE                       (RXSLIDE_MODE),                          

    //----------------------------------------------------------------------------------------------
    //  PCS Reserved Attributes
    //----------------------------------------------------------------------------------------------
    .PCS_RSVD0                          (PCS_RSVD0),
  
    //----------------------------------------------------------------------------------------------  
    //  PMA Reserved Attributes
    //----------------------------------------------------------------------------------------------      
    .TX_PMA_RSV0                        (16'h000A),                             
    .RX_PMA_RSV0                        (16'h00E0),                                        
      
    //----------------------------------------------------------------------------------------------
    //  CFOK Attributes                                                                 
    //----------------------------------------------------------------------------------------------              
    .RXCFOK_CFG0                        (16'b0011_1110_0000_0000),
    .RXCFOK_CFG1                        (16'b0000_0000_0100_0010),
    .RXCFOK_CFG2                        (16'b0000_0000_0010_1101),

    //----------------------------------------------------------------------------------------------
    //  RX CTLE
    //----------------------------------------------------------------------------------------------  
    .CTLE3_OCAP_EXT_CTRL	              ( 3'b000),                           
    .CTLE3_OCAP_EXT_EN	                ( 1'b0),                                
    .RX_EN_CTLE_RCAL_B                  ( 1'b0),                              

    //----------------------------------------------------------------------------------------------    
    //  RX LPM Attributes
    //----------------------------------------------------------------------------------------------        
    .RXLPM_CFG                          (16'b0000_0000_0000_0000),    
    .RXLPM_GC_CFG                       (16'b0000_0010_0000_0000),
    .RXLPM_KH_CFG0                      (16'b0000_0000_0000_0000),
    .RXLPM_KH_CFG1                      (16'b0000_0000_0000_0010),
    .RXLPM_OS_CFG0                      (16'b0000_0100_0000_0000),
    .RXLPM_OS_CFG1                      (16'b0000_0000_0000_0000),
 
    //----------------------------------------------------------------------------------------------    
    //  RX DFE Attributes
    //----------------------------------------------------------------------------------------------       
    .RXDFE_CFG0                         (16'b0100_1100_0000_0000), //(16'b0000110000000000),    [Changed for extracted model]
    .RXDFE_CFG1                         (16'b0000_0000_0000_0000),
    .RXDFE_GC_CFG0                      (16'b0001_1110_0000_0000), 
    .RXDFE_GC_CFG1                      (16'b0001_1001_0000_0000),  // different from GTH 
    .RXDFE_GC_CFG2                      (16'b0000_0000_0000_0000),  // different from GTH
    .RXDFE_H2_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_H2_CFG1                      (16'b0000_0000_0000_0010),
    .RXDFE_H3_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_H3_CFG1                      (16'b0000_0000_0000_0010),
    .RXDFE_H4_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_H4_CFG1                      (16'b0000_0000_0000_0011),
    .RXDFE_H5_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_H5_CFG1                      (16'b0000_0000_0000_0010),
    .RXDFE_H6_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_H6_CFG1                      (16'b0000_0000_0000_0010),
    .RXDFE_H7_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_H7_CFG1                      (16'b0000_0000_0000_0010), 
    .RXDFE_H8_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_H8_CFG1                      (16'b0000_0000_0000_0010),
    .RXDFE_H9_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_H9_CFG1                      (16'b0000_0000_0000_0010), 
    .RXDFE_HA_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_HA_CFG1                      (16'b0000_0000_0000_0010),
    .RXDFE_HB_CFG0                      (16'b0000_0000_0000_0000), //(16'b0010000000000000),    [Changed for extracted model]
    .RXDFE_HB_CFG1                      (16'b0000_0000_0000_0010),
    .RXDFE_HC_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_HC_CFG1                      (16'b0000_0000_0000_0010),
    .RXDFE_HD_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_HD_CFG1                      (16'b0000_0000_0000_0010),
    .RXDFE_HE_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_HE_CFG1                      (16'b0000_0000_0000_0010),
    .RXDFE_HF_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_HF_CFG1                      (16'b0000_0000_0000_0010),
    .RXDFE_OS_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_OS_CFG1                      (16'b0000_0000_0000_0010), //(16'b0000001000000000),    [Changed for extracted model]
    //.RXDFE_PWR_SAVING                   (16'b0),
    .RXDFE_UT_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_UT_CFG1                      (16'b0000_0000_0000_0010),
    .RXDFE_VP_CFG0                      (16'b0000_0000_0000_0000),
    .RXDFE_VP_CFG1                      (16'b0000_0000_0010_0010),
    .RXDFELPM_KL_CFG0                   (16'h0000),                  
    .RXDFELPM_KL_CFG1                   (16'h0022),             
    .RXDFELPM_KL_CFG2                   (16'h0100),                        
    //.RX_DFE_AGC_CFG0                    ( 2'b00),                               
    .RX_DFE_AGC_CFG1                    ( 2),  
    .RX_DFE_KL_LPM_KH_CFG0              ( 1),
    .RX_DFE_KL_LPM_KH_CFG1              ( 2),
    .RX_DFE_KL_LPM_KL_CFG0              ( 2'b01),
    .RX_DFE_KL_LPM_KL_CFG1              ( 3'b010),   
    .RX_DFELPM_CFG0                     ( 0),                                                            
    .RX_DFELPM_CFG1                     ( 1'b1),                                                               
    .RX_DFELPM_KLKH_AGC_STUP_EN         ( 1'b1),   
          
    //----------------------------------------------------------------------------------------------  
    //  TX PI attributes
    //----------------------------------------------------------------------------------------------
    .TX_PHICAL_CFG0	                    (16'h0000),                           
    .TX_PHICAL_CFG1	                    (16'h7e00),
    //.TX_PHICAL_CFG2	                    (16'h0000),
    .TX_PI_BIASSET	                    ( 0),                                  
    .TXPI_CFG0                          ( 2'b00),
    .TXPI_CFG1                          ( 2'b00),
    //.TXPI_CFG2                          ( 2'b00),
    //.TXPI_CFG3                          ( 1'b0),
    //.TXPI_CFG4                          ( 1'b1),
    //.TXPI_CFG5                          ( 3'b000),
    .TXPI_GRAY_SEL                      ( 1'b0),
    .TXPI_INVSTROBE_SEL                 ( 1'b0),
    //.TXPI_LPM                           ( 1'b0),
    .TXPI_PPM_CFG                       ( 8'b00000000),
    //.TXPI_PPMCLK_SEL                    ("TXUSRCLK2"),
    .TXPI_SYNFREQ_PPM                   ( 3'b000),
    //.TXPI_VREFSEL                       ( 1'b0),    
    
    //----------------------------------------------------------------------------------------------  
    //  RX PI Attributes
    //----------------------------------------------------------------------------------------------    
    //.RXPI_AUTO_BW_SEL_BYPASS            ( 1'b0),
    .RXPI_CFG0                          (16'h0100),
    .RXPI_CFG1                          (16'h0100),
    //.RXPI_LPM                           ( 1'b0),
    //.RXPI_SEL_LC                        ( 2'b00),
    //.RXPI_STARTCODE                     ( 2'b00),
    //.RXPI_VREFSEL                       ( 1'b0),              

    //----------------------------------------------------------------------------------------------
    //  RX CDR Attributes
    //----------------------------------------------------------------------------------------------    
    .CDR_SWAP_MODE_EN                   ( 1'b0),                 
    .RX_WIDEMODE_CDR                    ( 2'b01),                                      
    .RXCDR_CFG0                         (RXCDR_CFG0), 
    .RXCDR_CFG0_GEN3                    (RXCDR_CFG0_GEN3), 
    .RXCDR_CFG1                         (RXCDR_CFG1), 
    .RXCDR_CFG1_GEN3                    (RXCDR_CFG1_GEN3), 
    .RXCDR_CFG2                         (RXCDR_CFG2), 
    .RXCDR_CFG2_GEN3                    (RXCDR_CFG2_GEN3), 
    .RXCDR_CFG2_GEN4                    (RXCDR_CFG2_GEN4), 
    .RXCDR_CFG3                         (RXCDR_CFG3), 
    .RXCDR_CFG3_GEN3                    (RXCDR_CFG3_GEN3), 
    .RXCDR_CFG3_GEN4                    (RXCDR_CFG3_GEN4),
    .RXCDR_CFG4                         (RXCDR_CFG4), 
    .RXCDR_CFG4_GEN3                    (RXCDR_CFG4_GEN3), 
    .RXCDR_CFG5                         (RXCDR_CFG5), 
    .RXCDR_CFG5_GEN3                    (RXCDR_CFG5_GEN3), 
    .RXCDR_LOCK_CFG0                    (16'b1001_0000_1000_0001), 
    .RXCDR_LOCK_CFG1                    (16'b1001_0111_1110_0000), 
    .RXCDR_LOCK_CFG2                    (16'b0110_0100_0100_0001), 
    .RXCDR_LOCK_CFG3                    (16'b0000_0111_1110_0000), 

    //---------------------------------------------------------------------------------------------- 
    //  Eye Scan Attributes
    //----------------------------------------------------------------------------------------------
    .ES_CLK_PHASE_SEL                   ( 1'b0),                           
    .ES_CONTROL                         ( 6'b000000),                      
    .ES_ERRDET_EN                       ("FALSE"),                        
    .ES_EYE_SCAN_EN                     ("FALSE"),                        
    .ES_HORZ_OFFSET                     (12'b000000000000),                       
    .ES_PRESCALE                        ( 5'b00000),                                
    .ES_QUAL_MASK0                      (16'b0000000000000000),           
    .ES_QUAL_MASK1                      (16'b0000000000000000),           
    .ES_QUAL_MASK2                      (16'b0000000000000000),           
    .ES_QUAL_MASK3                      (16'b0000000000000000),           
    .ES_QUAL_MASK4                      (16'b0000000000000000),       
    .ES_QUAL_MASK5                      (16'b0000000000000000),           
    .ES_QUAL_MASK6                      (16'b0000000000000000),           
    .ES_QUAL_MASK7                      (16'b0000000000000000),           
    .ES_QUAL_MASK8                      (16'b0000000000000000),           
    .ES_QUAL_MASK9                      (16'b0000000000000000),         
    .ES_QUALIFIER0                      (16'b0000000000000000),           
    .ES_QUALIFIER1                      (16'b0000000000000000),           
    .ES_QUALIFIER2                      (16'b0000000000000000),           
    .ES_QUALIFIER3                      (16'b0000000000000000),           
    .ES_QUALIFIER4                      (16'b0000000000000000), 
    .ES_QUALIFIER5                      (16'b0000000000000000),           
    .ES_QUALIFIER6                      (16'b0000000000000000),           
    .ES_QUALIFIER7                      (16'b0000000000000000),           
    .ES_QUALIFIER8                      (16'b0000000000000000),           
    .ES_QUALIFIER9                      (16'b0000000000000000),   
    .ES_SDATA_MASK0                     (16'b0000000000000000),           
    .ES_SDATA_MASK1                     (16'b0000000000000000),           
    .ES_SDATA_MASK2                     (16'b0000000000000000),           
    .ES_SDATA_MASK3                     (16'b0000000000000000),           
    .ES_SDATA_MASK4                     (16'b0000000000000000), 
    .ES_SDATA_MASK5                     (16'b0000000000000000),           
    .ES_SDATA_MASK6                     (16'b0000000000000000),           
    .ES_SDATA_MASK7                     (16'b0000000000000000),           
    .ES_SDATA_MASK8                     (16'b0000000000000000),   
    .ES_SDATA_MASK9                     (16'b0000000000000000),          
    .EYE_SCAN_SWAP_EN                   ( 1'b0),
    .RX_EYESCAN_VS_CODE                 ( 7'b0000000),
    .RX_EYESCAN_VS_NEG_DIR              ( 1'b0),
    .RX_EYESCAN_VS_RANGE                ( 2'b00),
    .RX_EYESCAN_VS_UT_SIGN              ( 1'b0),                        
  
    //----------------------------------------------------------------------------------------------
    //  Loopback & PRBS Attributes
    //----------------------------------------------------------------------------------------------
    .RXPRBS_ERR_LOOPBACK                ( 1'b0),     
    .RXPRBS_LINKACQ_CNT                 (15),                                                   
                                                                                                    
    //----------------------------------------------------------------------------------------------   
    //  Digital Monitor Attribute
    //----------------------------------------------------------------------------------------------                     
    .DMONITOR_CFG0                      (10'b0000000000),                                                  
    .DMONITOR_CFG1                      ( 8'b00000000),                                                   
                                                      
    //----------------------------------------------------------------------------------------------   
    //  AC JTAG Attributes
    //----------------------------------------------------------------------------------------------                     
    .ACJTAG_DEBUG_MODE                  ( 1'b0),                                                        
    .ACJTAG_MODE                        ( 1'b0),                                                        
    .ACJTAG_RESET                       ( 1'b0),      
    
    //----------------------------------------------------------------------------------------------
    //  USB Attributes
    //----------------------------------------------------------------------------------------------                 
    .USB_BOTH_BURST_IDLE                ( 1'b0),
    .USB_BURSTMAX_U3WAKE	              ( 7'b1111111),
    .USB_BURSTMIN_U3WAKE	              ( 7'b1100011),
    .USB_CLK_COR_EQ_EN                  ( 1'b1),                              
    .USB_EXT_CNTL                       ( 1'b1),
    .USB_IDLEMAX_POLLING                (10'b1010111011),
    .USB_IDLEMIN_POLLING                (10'b0100101011),
    .USB_LFPS_TPERIOD	                  ( 4'b0011),
    .USB_LFPS_TPERIOD_ACCURATE	        ( 1'b1),
    .USB_LFPSPING_BURST	                ( 9'b000000101),
    .USB_LFPSPOLLING_BURST	            ( 9'b000110001),
    .USB_LFPSPOLLING_IDLE_MS	          ( 9'b000000100),
    .USB_LFPSU1EXIT_BURST	              ( 9'b000011101),
    .USB_LFPSU2LPEXIT_BURST_MS	        ( 9'b001100011),
    .USB_LFPSU3WAKE_BURST_MS	          ( 9'b111110011),
    .USB_MODE                           (USB_MODE), 
    .USB_PCIE_ERR_REP_DIS               ( 1'b0),                                // For Debug
    .USB_PING_SATA_MAX_INIT             (21),
    .USB_PING_SATA_MIN_INIT             (12),
    .USB_POLL_SATA_MAX_BURST            ( 8),
    .USB_POLL_SATA_MIN_BURST            ( 4),
    .USB_RAW_ELEC                       ( 1'b1),                               
    .USB_RXIDLE_P0_CTRL                 ( 1'b1),
    .USB_TXIDLE_TUNE_ENABLE             ( 1'b1),
    .USB_U1_SATA_MAX_WAKE               ( 7),
    .USB_U1_SATA_MIN_WAKE               ( 4),
    .USB_U2_SAS_MAX_COM                 (64),   
    .USB_U2_SAS_MIN_COM                 (36),
    
    //---------------------------------------------------------------------------------------------- 
    //  SAS & SATA Attributes (Not used)
    //---------------------------------------------------------------------------------------------- 
  //.SAS12G_MODE                        ( 1'b0),
  //.SATA_BURST_SEQ_LEN                 ( 4'b1111),
  //.SATA_BURST_VAL                     ( 3'b100),
  //.SATA_CPLL_CFG                      ("VCO_3000MHZ"),
  //.SATA_EIDLE_VAL                     ( 3'b100), 
            
    //---------------------------------------------------------------------------------------------- 
    //  CKCAL Attributes
    //---------------------------------------------------------------------------------------------- 
    .CKCAL1_CFG_0	                      (16'hC0C0), //(16'b0000000000000000), [Changed for extracted model]
    .CKCAL1_CFG_1	                      (16'h00C0), //(16'b0000000000000000), [Changed for extracted model] 
    .CKCAL1_CFG_2	                      (16'b0000000000000000),
    .CKCAL1_CFG_3	                      (16'b0000000000000000),
    .CKCAL2_CFG_0	                      (16'h8181), //(16'b0000000000000000), [Changed for extracted model]
    .CKCAL2_CFG_1	                      (16'h8081), //(16'b0000000000000000), [Changed for extracted model]
    .CKCAL2_CFG_2	                      (16'b0000000000000000),
    .CKCAL2_CFG_3	                      (16'b0000000000000000),
    .CKCAL2_CFG_4	                      (16'b0000000000000000),
    //.CKCAL_RSVD0	                      (16'h4000),
    //.CKCAL_RSVD1	                      (16'h0000),
    .RXCKCAL1_I_LOOP_RST_CFG	          (16'h0000),
    .RXCKCAL1_IQ_LOOP_RST_CFG	          (16'h0000),
    .RXCKCAL1_Q_LOOP_RST_CFG	          (16'h0000),
    .RXCKCAL2_D_LOOP_RST_CFG	          (16'h0000),
    .RXCKCAL2_DX_LOOP_RST_CFG	          (16'h0000),
    .RXCKCAL2_S_LOOP_RST_CFG	          (16'h0000),
    .RXCKCAL2_X_LOOP_RST_CFG	          (16'h0000),
  
    //----------------------------------------------------------------------------------------------
    //  Summer Attributes
    //----------------------------------------------------------------------------------------------
    .RX_SUM_DFETAPREP_EN                ( 1'b0),
    .RX_SUM_IREF_TUNE                   ( 4'b0000),
    .RX_SUM_VCM_OVWR                    ( 1'b0),
    .RX_SUM_VCMTUNE                     ( 4'b1000),
    .RX_SUM_VREF_TUNE                   ( 3'b100),

    //----------------------------------------------------------------------------------------------
    //  Attributes
    //----------------------------------------------------------------------------------------------                 
    .A_RXOSCALRESET                     ( 1'b0),   
    .A_RXPROGDIVRESET                   ( 1'b0),
    .A_RXTERMINATION                    ( 1'b1),
    .A_TXDIFFCTRL                       ( 5'b11111),
    .A_TXPROGDIVRESET                   ( 1'b0),
    .ADAPT_CFG0                         ( 16'b1001001000000000),
    .ADAPT_CFG1                         ( 16'b1000000000011100),
    .ADAPT_CFG2                         ( 16'b0000000000000000), 
    //.CAPBYPASS_FORCE                    ( 1'b0),                                
    .CH_HSPMUX                          ( 16'h0000),
    .DDI_CTRL                           ( 2'b00),
    .DDI_REALIGN_WAIT                   (15),
    .DELAY_ELEC                         ( 1'b0),                              
    .ISCAN_CK_PH_SEL2                   ( 1'b0),                                
    .PREIQ_FREQ_BST                     ( 0),                                   
    //.PROCESS_PAR                        ( 3'b010), 
    .RX_CAPFF_SARC_ENB                  ( 1'b0),    
    .RX_DDI_SEL                         ( 6'b000000),  
    .RX_DEGEN_CTRL                      ( 3'b011),                              
    //.RX_DIV2_MODE_B                     ( 1'b0),                                
    //.RX_EN_HI_LR                        ( 1'b0),
    //.RX_EXT_RL_CTRL                     ( 9'b000000000),                        
    .RX_RESLOAD_CTRL	                  ( 4'b0000),                             
    .RX_RESLOAD_OVRD	                  ( 1'b0),                                
    .RX_VREG_CTRL	                      ( 3'b101),                              
    .RX_VREG_PDB	                      ( 1'b1),                                
    .RX_XMODE_SEL	                      ( 1'b0),                                
    .TAPDLY_SET_TX                      ( 2'b00),
    //.TEMPERATURE_PAR                    ( 4'b0010),
    .TST_RSV0                           ( 8'b00000000),                                     
    .TST_RSV1                           ( 8'b00000000),
    .TX_DCC_LOOP_RST_CFG                (16'h0000),                             
    //.TX_DRVMUX_CTRL                     ( 2),                                   
    //.TX_PREDRV_CTRL                     ( 2),                                   
    .TX_PMADATA_OPT                     ( 1'b0)    
)                                                                                                   
gtye4_channel_smsw_i                                                                                     
(                                                                                                                                                                                                   
    //----------------------------------------------------------------------------------------------
    //  Clock Ports
    //----------------------------------------------------------------------------------------------
    .GTGREFCLK                          ( 1'd0),                                                     
    .GTREFCLK0                          (GT_GTREFCLK0),                                            
    .GTREFCLK1                          ( 1'd0),                                                    
    .GTNORTHREFCLK0                     ( 1'd0),                                                    
    .GTNORTHREFCLK1                     ( 1'd0),                                                    
    .GTSOUTHREFCLK0                     ( 1'd0),                                                    
    .GTSOUTHREFCLK1                     ( 1'd0),                                             
    .TXUSRCLK                           (GT_TXUSRCLK),                                              
    .RXUSRCLK                           (GT_RXUSRCLK),                                              
    .TXUSRCLK2                          (GT_TXUSRCLK2),                                             
    .RXUSRCLK2                          (GT_RXUSRCLK2),  
    .TXPLLCLKSEL                        (PLLCLKSEL),            
    .RXPLLCLKSEL                        (PLLCLKSEL),                                                    
    .TXSYSCLKSEL                        (SYSCLKSEL),                                             
    .RXSYSCLKSEL                        (SYSCLKSEL),                             
    .TXOUTCLKSEL                        (GT_TXOUTCLKSEL), //( 3'd5),            // Select TXPROGDIVCLK
    .RXOUTCLKSEL                        ( 3'd2),                                // Select RXOUTCLKPMA
    .CLKRSVD0                           ( 1'd0),          
    .CLKRSVD1                           ( 1'd0),            
                                                                                                   
    .TXOUTCLK                           (GT_TXOUTCLK),                                             
    .RXOUTCLK                           (GT_RXOUTCLK),                                                        
    .TXOUTCLKFABRIC                     (GT_TXOUTCLKFABRIC),                                                        
    .RXOUTCLKFABRIC                     (GT_RXOUTCLKFABRIC),                                                        
    .TXOUTCLKPCS                        (GT_TXOUTCLKPCS),                                                        
    .RXOUTCLKPCS                        (GT_RXOUTCLKPCS),  
    .RXRECCLKOUT                        (GT_RXRECCLKOUT),                                                    
    .GTREFCLKMONITOR                    (),                                 
    
    //----------------------------------------------------------------------------------------------
    //  BUFG_GT Controller Ports
    //----------------------------------------------------------------------------------------------
    .BUFGTCE                            (GT_BUFGTCE),      
    .BUFGTCEMASK                        (GT_BUFGTCEMASK), 
    .BUFGTDIV                           (GT_BUFGTDIV), 
    .BUFGTRESET                         (GT_BUFGTRESET), 
    .BUFGTRSTMASK                       (GT_BUFGTRSTMASK),       
    
    //----------------------------------------------------------------------------------------------
    //  CPLL Ports
    //----------------------------------------------------------------------------------------------
    .CPLLFREQLOCK                       (GT_MASTER_CPLLLOCK),                 
    .CPLLLOCKDETCLK                     ( 1'd0),                              
    .CPLLLOCKEN                         ( 1'd1),    
    .CPLLPD                             (GT_CPLLPD),    
    .CPLLREFCLKSEL                      ( 3'd1),                               
    .CPLLRESET                          (GT_CPLLRESET),                               
  
    .CPLLFBCLKLOST                      (),     
    .CPLLLOCK                           (GT_CPLLLOCK),                                            
    .CPLLREFCLKLOST                     (),                    
             
    //----------------------------------------------------------------------------------------------
    //  QPLL Ports                                                                                   
    //----------------------------------------------------------------------------------------------
    .QPLL0CLK                           (GT_QPLL0CLK),                           
    .QPLL0REFCLK                        (GT_QPLL0REFCLK),                        
    .QPLL0FREQLOCK                      (GT_QPLL0LOCK),                         
    .QPLL1CLK                           (GT_QPLL1CLK),  
    .QPLL1REFCLK                        (GT_QPLL1REFCLK),           
    .QPLL1FREQLOCK                      (GT_QPLL1LOCK),                         
    
    //----------------------------------------------------------------------------------------------
    //  Reset Ports
    //----------------------------------------------------------------------------------------------                                                                                                                             
    .GTTXRESET                          (GT_GTTXRESET),                                             
    .GTRXRESET                          (GT_GTRXRESET),  
    .GTRXRESETSEL                       ( 1'd0),                                
    .GTTXRESETSEL                       ( 1'd0),                                
    .TXPROGDIVRESET                     (GT_TXPROGDIVRESET),                       
    .RXPROGDIVRESET                     ( 1'd0),                                                                            
    .TXPMARESET                         (GT_TXPMARESET),                                            
    .RXPMARESET                         (GT_RXPMARESET),                                            
    .TXPCSRESET                         (GT_TXPCSRESET),   
    .RXPCSRESET                         (GT_RXPCSRESET),   
    .TXUSERRDY                          (GT_TXUSERRDY),                                             
    .RXUSERRDY                          (GT_RXUSERRDY),   
    .CFGRESET                           ( 1'd0),                                                    
    .RESETOVRD                          ( GT_RESETOVRD),  
    .RXOOBRESET                         ( 1'd0),                                              
                                           
    .GTPOWERGOOD                        (GT_GTPOWERGOOD), 
    .TXPRGDIVRESETDONE                  (GT_TXPROGDIVRESETDONE),
    .RXPRGDIVRESETDONE                  (),        
    .TXPMARESETDONE                     (GT_TXPMARESETDONE),    
    .RXPMARESETDONE                     (GT_RXPMARESETDONE),                                                                                                      
    .TXRESETDONE                        (GT_TXRESETDONE),                                           
    .RXRESETDONE                        (GT_RXRESETDONE),  
    .RESETEXCEPTION                     (),

    //----------------------------------------------------------------------------------------------
    //  PCIe Ports
    //----------------------------------------------------------------------------------------------
    .PCIERSTIDLE                        (GT_PCIERSTIDLE),        
    .PCIERSTTXSYNCSTART                 (GT_PCIERSTTXSYNCSTART), 
    .PCIEEQRXEQADAPTDONE                (GT_PCIEEQRXEQADAPTDONE),
    .PCIEUSERRATEDONE                   (GT_PCIEUSERRATEDONE),
             
    .PCIEUSERPHYSTATUSRST               (GT_PCIEUSERPHYSTATUSRST),    
    .PCIERATEQPLLPD                     (GT_PCIERATEQPLLPD),                    
    .PCIERATEQPLLRESET                  (GT_PCIERATEQPLLRESET),                 
    .PCIERATEIDLE                       (GT_PCIERATEIDLE),            
    .PCIESYNCTXSYNCDONE                 (GT_PCIESYNCTXSYNCDONE),                          
    .PCIERATEGEN3                       (pcierategen3),    
    .PCIEUSERGEN3RDY                    (GT_PCIEUSERGEN3RDY),   
    .PCIEUSERRATESTART                  (GT_PCIEUSERRATESTART),    
           
    //----------------------------------------------------------------------------------------------
    //  Serial Line Ports
    //----------------------------------------------------------------------------------------------
    .GTYRXP                             (GT_RXP),                                                   
    .GTYRXN                             (GT_RXN),   
   
    .GTYTXP                             (GT_TXP),                                                 
    .GTYTXN                             (GT_TXN),   

    //----------------------------------------------------------------------------------------------
    //  TX Data Ports
    //----------------------------------------------------------------------------------------------
    .TXDATA                             (txdata),                                     
    .TXCTRL0                            (txctrl0),
    .TXCTRL1                            (txctrl1),  
    .TXCTRL2                            (txctrl2),
    .TXDATAEXTENDRSVD                   ( 8'd0),                                

    //----------------------------------------------------------------------------------------------
    //  RX Data Ports
    //----------------------------------------------------------------------------------------------
    .RXDATA                             (rxdata),                                                    
    .RXCTRL0                            (rxctrl0),   
    .RXCTRL1                            (), 
    .RXCTRL2                            (),
    .RXCTRL3                            (), 
    .RXDATAEXTENDRSVD                   (),                                     
 
    //----------------------------------------------------------------------------------------------
    //  PHY Command Ports
    //----------------------------------------------------------------------------------------------
    .TXDETECTRX                         (GT_TXDETECTRX),                                            
    .TXELECIDLE                         (GT_TXELECIDLE),                                      
    .TXPDELECIDLEMODE                   ( 1'd0),                                                                                 
    .RXELECIDLEMODE                     ( 2'd0),                                
    .SIGVALIDCLK                        ( 1'd0),                                                                                    
    .TXPOLARITY                         ( 1'd0),                                              
    .RXPOLARITY                         (GT_RXPOLARITY),                                
    .TXPD                               (GT_POWERDOWN),                                           
    .RXPD                               (GT_POWERDOWN),                                           
    .TXRATE                             ({1'd0, GT_RATE}),                                                
    .RXRATE                             ({1'd0, GT_RATE}),                                                
    .TXRATEMODE                         ( 1'd0),                                                    
    .RXRATEMODE                         ( 1'd0),                                                    
 
    //----------------------------------------------------------------------------------------------
    //  PHY Status Ports
    //----------------------------------------------------------------------------------------------
    .RXVALID                            (GT_RXVALID),                                              
    .PHYSTATUS                          (GT_PHYSTATUS),                                            
    .RXELECIDLE                         (rxelecidle_int),                                           
    .RXSTATUS                           (GT_RXSTATUS),                                             
    .TXRATEDONE                         (),                                           
    .RXRATEDONE                         (GT_RXRATEDONE),                  
 
    //----------------------------------------------------------------------------------------------
    //  TX Driver Ports
    //----------------------------------------------------------------------------------------------
    .TXMARGIN                           (GT_TXMARGIN),                                           
    .TXSWING                            (GT_TXSWING),                                            
    .TXDEEMPH                           (GT_TXDEEMPH),                                                                     
    .TXDIFFCTRL                         ( 5'b11111),
    .TXINHIBIT                          ( 1'd0),                                                  

    //----------------------------------------------------------------------------------------------
    //  TX Driver Ports (Gen3)
    //----------------------------------------------------------------------------------------------
    .TXPRECURSOR                        (GT_TXPRECURSOR),                                          
    .TXMAINCURSOR                       (GT_TXMAINCURSOR),                                         
    .TXPOSTCURSOR                       (GT_TXPOSTCURSOR),                                                                                     

    //----------------------------------------------------------------------------------------------
    //  PCS Reserved Ports
    //---------------------------------------------------------------------------------------------- 
    .PCSRSVDIN                          (16'h0001),                             // CHECK                                                                               
    .PCSRSVDOUT                         (pcsrsvdout),     
    
    //----------------------------------------------------------------------------------------------
    //  RX Monitor Ports
    //----------------------------------------------------------------------------------------------
    .RXMONITORSEL                       ( 2'd0), 
    .RXMONITOROUT                       (),                                                                                                                                                                                                            
                                                                 
    //----------------------------------------------------------------------------------------------
    //  Comma Detect & Align Ports
    //----------------------------------------------------------------------------------------------
    .RXCOMMADETEN                       ( 1'd1),                  
    .RXMCOMMAALIGNEN                    (!pcierategen3),          
    .RXPCOMMAALIGNEN                    (!pcierategen3),          
                                                                                 
    .RXCOMMADET                         (),                                            
    .RXBYTEISALIGNED                    (),                                        
    .RXBYTEREALIGN                      (),                                                                                                                 
                                                                                                    
    //----------------------------------------------------------------------------------------------
    // 8B10B Ports
    //----------------------------------------------------------------------------------------------
    .TX8B10BBYPASS                      ( 8'd0),                                                  
    .TX8B10BEN                          (!pcierategen3),                            
    .RX8B10BEN                          (!pcierategen3),                            
           
    //----------------------------------------------------------------------------------------------
    //  TX Buffer Ports
    //----------------------------------------------------------------------------------------------
    .TXBUFSTATUS                        (),                                                        
                                                                                                    
    //----------------------------------------------------------------------------------------------
    //  RX Buffer Ports
    //----------------------------------------------------------------------------------------------
    .RXBUFRESET                         (GT_RXBUFRESET),                                          
    .RXBUFSTATUS                        (),                
                      
    //----------------------------------------------------------------------------------------------
    //  Clock Correction Ports
    //----------------------------------------------------------------------------------------------
    .RXCLKCORCNT                        (),                            
                    
    //----------------------------------------------------------------------------------------------
    //  Channel Bonding Ports (disable)
    //----------------------------------------------------------------------------------------------
    .RXCHBONDEN                         ( 1'd0),                                         
    .RXCHBONDI                          ( 5'd0),                                         
    .RXCHBONDLEVEL                      ( 3'd0),                                         
    .RXCHBONDMASTER                     ( 1'd0),                                         
    .RXCHBONDSLAVE                      ( 1'd0),                                         
                                                                                    
    .RXCHANBONDSEQ                      (),                                         
    .RXCHANISALIGNED                    (),                                         
    .RXCHANREALIGN                      (),                                         
    .RXCHBONDO                          (),                                                                                                                                                                       
 
    //----------------------------------------------------------------------------------------------
    //  TX Phase Alignment Ports
    //----------------------------------------------------------------------------------------------
    .TXPHALIGN                          ( 1'd0),
    .TXPHALIGNEN                        ( 1'd0),
    .TXPHDLYPD                          ( 1'd0),
    .TXPHDLYRESET                       ( 1'd0),
    .TXPHDLYTSTCLK                      ( 1'd0),
    .TXPHINIT                           ( 1'd0),
    .TXPHOVRDEN                         ( 1'd0),
   
    .TXPHALIGNDONE                      (GT_TXPHALIGNDONE),
    .TXPHINITDONE                       (),
   
    //----------------------------------------------------------------------------------------------
    //  TX Delay Alignment Ports
    //----------------------------------------------------------------------------------------------
    .TXDLYBYPASS                        ( 1'd0),
    .TXDLYEN                            ( 1'd0),
    .TXDLYHOLD                          ( 1'd0),
    .TXDLYOVRDEN                        ( 1'd0),
    .TXDLYSRESET                        ( 1'd0),
    .TXDLYUPDOWN                        ( 1'd0),
       
    .TXDLYSRESETDONE                    (),       
          
    //----------------------------------------------------------------------------------------------
    //  TX Auto Sync Alignment Ports 
    //----------------------------------------------------------------------------------------------
    .TXSYNCALLIN                        (GT_TXSYNCALLIN),
    .TXSYNCIN                           (GT_TXSYNCIN),
    .TXSYNCMODE                         (MASTER_LANE),                                         
                
    .TXSYNCDONE                         (),
    .TXSYNCOUT                          (GT_TXSYNCOUT),

    //----------------------------------------------------------------------------------------------
    //  RX Phase Alignment Ports (disable)
    //----------------------------------------------------------------------------------------------
    .RXPHALIGN                          ( 1'd0),
    .RXPHALIGNEN                        ( 1'd0),
    .RXPHDLYPD                          ( 1'd0),
    .RXPHDLYRESET                       ( 1'd0),
  //.RXPHOVRDEN                         ( 1'd0),
   
    .RXPHALIGNDONE                      (),
    .RXPHALIGNERR                       (),
       
    //----------------------------------------------------------------------------------------------
    //  RX Delay Alignment Ports (disable)
    //----------------------------------------------------------------------------------------------
    .RXDLYBYPASS                        ( 1'd1),
    .RXDLYEN                            ( 1'd0),
    .RXDLYOVRDEN                        ( 1'd0),
    .RXDLYSRESET                        ( 1'd0),
   
    .RXDLYSRESETDONE                    (),                                           
        
    //----------------------------------------------------------------------------------------------
    //  RX Auto Sync Alignment Ports (disable)
    //----------------------------------------------------------------------------------------------
    .RXSYNCALLIN                        ( 1'd0),
    .RXSYNCIN                           ( 1'd0),
    .RXSYNCMODE                         ( 1'd0),                                                    
                                                                                                    
    .RXSYNCDONE                         (),                                                
    .RXSYNCOUT                          (),    
       
    //----------------------------------------------------------------------------------------------
    //  Gearbox Ports 
    //----------------------------------------------------------------------------------------------
    .TXHEADER                           ( 6'd0), 
    .TXLATCLK                           ( 1'd0),                                                    
    .TXSEQUENCE                         ( 7'd0),                                                    
    .RXGEARBOXSLIP                      ( 1'd0),  
    .RXLATCLK                           ( 1'd0),  
    .RXSLIDE                            ( 1'd0),                                                    
                                                                                                    
    .RXDATAVALID                        (),                 
    .RXHEADER                           (),                                                         
    .RXHEADERVALID                      (), 
    .RXSLIDERDY                         (),                                                         
    .RXSTARTOFSEQ                       (),                             
                   
    //----------------------------------------------------------------------------------------------
    //  RX Slip Ports 
    //----------------------------------------------------------------------------------------------
    .RXSLIPOUTCLK                       ( 1'd0),
    .RXSLIPPMA                          ( 1'd0),   
                                                                   
    .RXSLIPDONE                         (),     
    .RXSLIPOUTCLKRDY                    (),
    .RXSLIPPMARDY                       (),             
       
    //----------------------------------------------------------------------------------------------
    //  RX LPM Ports 
    //----------------------------------------------------------------------------------------------
    .RXLPMEN                            (!pcierategen3),    
    .RXLPMGCHOLD                        ( 1'b0),            
    .RXLPMGCOVRDEN                      ( 1'b0),
    .RXLPMHFHOLD                        ( 1'b0),            
    .RXLPMHFOVRDEN                      ( 1'b0),
    .RXLPMLFHOLD                        ( 1'b0),         
    .RXLPMLFKLOVRDEN                    ( 1'b0), 
    .RXLPMOSHOLD                        ( 1'b0),            
    .RXLPMOSOVRDEN                      ( 1'b0),
                                                                                                    
    //----------------------------------------------------------------------------------------------
    //  RX DFE Ports
    //----------------------------------------------------------------------------------------------
    ////.RXDFEAGCCTRL                       ( 2'h1), //( 2'b00),     [Changed for extracted model]
    .RXDFEAGCHOLD                       ( 1'b0),            
    .RXDFEAGCOVRDEN                     ( 1'b0),
    .RXDFECFOKFCNUM                     ( 4'b0000),                             
    .RXDFECFOKFEN                       ( 1'b0),                                
    .RXDFECFOKFPULSE                    ( 1'b0),                                
    .RXDFECFOKHOLD                      ( 1'b0),                                
    .RXDFECFOKOVREN                     ( 1'b0),                                
    .RXDFEKHHOLD                        ( 1'b0),
    .RXDFEKHOVRDEN                      ( 1'b0),
    .RXDFELFHOLD                        ( 1'b0),          
    .RXDFELFOVRDEN                      ( 1'b0),
    .RXDFELPMRESET                      (GT_RXDFELPMRESET),
    .RXDFETAP2HOLD                      ( 1'b0),
    .RXDFETAP2OVRDEN                    ( 1'b0),
    .RXDFETAP3HOLD                      ( 1'b0),
    .RXDFETAP3OVRDEN                    ( 1'b0),
    .RXDFETAP4HOLD                      ( 1'b0),
    .RXDFETAP4OVRDEN                    ( 1'b0),
    .RXDFETAP5HOLD                      ( 1'b0),
    .RXDFETAP5OVRDEN                    ( 1'b0),
    .RXDFETAP6HOLD                      ( 1'b0),
    .RXDFETAP6OVRDEN                    ( 1'b0),
    .RXDFETAP7HOLD                      ( 1'b0),
    .RXDFETAP7OVRDEN                    ( 1'b0),
    .RXDFETAP8HOLD                      ( 1'b0),
    .RXDFETAP8OVRDEN                    ( 1'b0),
    .RXDFETAP9HOLD                      ( 1'b0),
    .RXDFETAP9OVRDEN                    ( 1'b0),
    .RXDFETAP10HOLD                     ( 1'b0),
    .RXDFETAP10OVRDEN                   ( 1'b0),
    .RXDFETAP11HOLD                     ( 1'b0),
    .RXDFETAP11OVRDEN                   ( 1'b0),
    .RXDFETAP12HOLD                     ( 1'b0),
    .RXDFETAP12OVRDEN                   ( 1'b0),
    .RXDFETAP13HOLD                     ( 1'b0),
    .RXDFETAP13OVRDEN                   ( 1'b0),
    .RXDFETAP14HOLD                     ( 1'b0),
    .RXDFETAP14OVRDEN                   ( 1'b0),
    .RXDFETAP15HOLD                     ( 1'b0),
    .RXDFETAP15OVRDEN                   ( 1'b0),
    .RXDFEUTHOLD                        ( 1'b0),
    .RXDFEUTOVRDEN                      ( 1'b0),
    .RXDFEVPHOLD                        ( 1'b0),
    .RXDFEVPOVRDEN                      ( 1'b0),
    .RXDFEXYDEN                         ( 1'b1),                                                                                                    
    
    //----------------------------------------------------------------------------------------------
    //  TX PI Ports
    //----------------------------------------------------------------------------------------------
    .TXPIPPMEN                          ( 1'd0),
    .TXPIPPMOVRDEN                      ( 1'd0),
    .TXPIPPMPD                          ( 1'd0),
    .TXPIPPMSEL                         ( 1'd0),
    .TXPIPPMSTEPSIZE                    ( 5'd0),
    .TXPISOPD                           ( 1'd0),   
    
    //----------------------------------------------------------------------------------------------
    //  RX CDR Ports
    //----------------------------------------------------------------------------------------------
    .CDRSTEPDIR                         ( 1'b0),                                 
    .CDRSTEPSQ                          ( 1'b0),                                
    .CDRSTEPSX                          ( 1'b0),                               
    .RXCDRFREQRESET                     (GT_RXCDRFREQRESET),
    .RXCDRHOLD                          (GT_RXCDRHOLD),
    .RXCDROVRDEN                        ( 1'd0),
    .RXCDRRESET                         (rxcdrreset_int),
    
    .RXCDRLOCK                          (GT_RXCDRLOCK),    
    .RXCDRPHDONE                        (), 
       
    //----------------------------------------------------------------------------------------------
    //  Eye Scan Ports
    //----------------------------------------------------------------------------------------------                                          
    .EYESCANRESET                       ( 1'd0),                                             
    .EYESCANTRIGGER                     ( 1'd0),                                             
                                                                                            
    .EYESCANDATAERROR                   (),           
       
    //----------------------------------------------------------------------------------------------
    //  RX OS Ports
    //----------------------------------------------------------------------------------------------
    .RXOSCALRESET                       ( 1'b0),
    .RXOSHOLD                           ( 1'b0),
    .RXOSOVRDEN                         ( 1'b0),    
 
    .RXOSINTDONE                        (),                                                         
    .RXOSINTSTARTED                     (),                                                         
    .RXOSINTSTROBEDONE                  (),                                                         
    .RXOSINTSTROBESTARTED               (),         
           
    //----------------------------------------------------------------------------------------------
    //  DRP Ports
    //----------------------------------------------------------------------------------------------
    .DRPCLK                             (GT_DRPCLK), 
    .DRPRST                             ( 1'd0),                                                                                
    .DRPADDR                            (GT_DRPADDR),                                                    
    .DRPEN                              (GT_DRPEN),                                                    
    .DRPWE                              (GT_DRPWE), 
    .DRPDI                              (GT_DRPDI),                                                    
        
    .DRPRDY                             (GT_DRPRDY),                                                         
    .DRPDO                              (GT_DRPDO),

    //----------------------------------------------------------------------------------------------
    //  Loopback & PRBS Ports
    //----------------------------------------------------------------------------------------------
    .LOOPBACK                           (GT_LOOPBACK),      
    .TXPRBSSEL                          (GT_PRBSSEL),                                                    
    .RXPRBSSEL                          (GT_PRBSSEL),  
    .TXPRBSFORCEERR                     (GT_TXPRBSFORCEERR),  
    .RXPRBSCNTRESET                     (GT_RXPRBSCNTRESET),  
                   
    .RXPRBSERR                          (GT_RXPRBSERR),                                                
    .RXPRBSLOCKED                       (GT_RXPRBSLOCKED),       

    //----------------------------------------------------------------------------------------------
    //  Digital Monitor Ports                                                                             
    //----------------------------------------------------------------------------------------------
    .DMONFIFORESET                      ( 1'd0),                                                    
    .DMONITORCLK                        ( 1'd0),                                                    
    
    .DMONITOROUT                        (),    
    .DMONITOROUTCLK                     (),                                             
      
    //----------------------------------------------------------------------------------------------
    //  USB Ports
    //----------------------------------------------------------------------------------------------
    .TXONESZEROS                        (GT_TXONESZEROS),
    .RXEQTRAINING                       (GT_RXEQTRAINING),
    .RXTERMINATION                      (GT_RXTERMINATION),    
    
    .POWERPRESENT                       (GT_POWERPRESENT),           
        
    //----------------------------------------------------------------------------------------------
    //  USB LFPS Ports
    //----------------------------------------------------------------------------------------------
    .TXLFPSTRESET                       ( 1'b0),      
    .TXLFPSU2LPEXIT                     ( 1'b0),
    .TXLFPSU3WAKE                       ( 1'b0),
    
    .RXLFPSTRESETDET                    (),             
    .RXLFPSU2LPEXITDET                  (),             
    .RXLFPSU3WAKEDET                    (),            
      
    //----------------------------------------------------------------------------------------------
    //  SATA Ports 
    //----------------------------------------------------------------------------------------------
    .TXCOMINIT                          ( 1'd0),                                                    
    .TXCOMSAS                           ( 1'd0),                                                    
    .TXCOMWAKE                          ( 1'd0),                                                    

    .TXCOMFINISH                        (),                                                         
    .RXCOMINITDET                       (),                                                         
    .RXCOMSASDET                        (),                                                         
    .RXCOMWAKEDET                       (),                                                    

    //----------------------------------------------------------------------------------------------
    //  QPI
    //----------------------------------------------------------------------------------------------
    ////.RXQPIEN                            ( 1'd0),
    ////.TXQPIBIASEN                        ( 1'b0),                                
    ////.TXQPIWEAKPUP                       ( 1'b0),                              
    
    ////.RXQPISENN                          (),
    ////.RXQPISENP                          (),
    ////.TXQPISENN                          (),
    ////.TXQPISENP                          (),

    //----------------------------------------------------------------------------------------------
    //  GT Ports
    //----------------------------------------------------------------------------------------------
    .FREQOS                             ( 1'd0),    
    .GTRSVD                             (16'd0),
    .INCPCTRL                           ( 1'd0),
    .RXAFECFOKEN                        ( 1'd0),                                
    .RXCKCALRESET                       ( 1'b0),                                
    .RXCKCALSTART                       ( 7'd0),                                
    .TSTIN                              (20'h00000),                                                
    .TXDCCFORCESTART                    ( 1'b0),                                
    .TXDCCRESET                         ( 1'b0),                                
    .TXMUXDCDEXHOLD                     ( 1'b0),                                
    .TXMUXDCDORWREN                     ( 1'b0),                                
                                                                                   
    .PINRSRVDAS                         (),                                     
    .RXCKCALDONE                        (),                                     
    .TXDCCDONE                          ()                                      
);

end else begin: GTH_CHANNEL
//--------------------------------------------------------------------------------------------------
//  GTH Channel
//--------------------------------------------------------------------------------------------------
GTHE4_CHANNEL #
(  
    //----------------------------------------------------------------------------------------------
    //  Simulation Attributes
    //----------------------------------------------------------------------------------------------
    .SIM_MODE                           ("FAST"),                                    
    .SIM_RECEIVER_DETECT_PASS           ("TRUE"),
    .SIM_RESET_SPEEDUP                  ("TRUE"),
    .SIM_TX_EIDLE_DRIVE_LEVEL           (SIM_TX_EIDLE_DRIVE_LEVEL),
  //.SIM_VERSION                        (1),                             
   
    //----------------------------------------------------------------------------------------------     
    //  Clock Attributes
    //----------------------------------------------------------------------------------------------                       
    .TXREFCLKDIV2_SEL                   ( 1'b0),                              
    .RXREFCLKDIV2_SEL                   ( 1'b0),                                
    .TX_CLK25_DIV                       (CLK25_DIV),                                                    
    .RX_CLK25_DIV                       (CLK25_DIV),                                                    
    .TX_CLKMUX_EN                       ( 1'b1),                                                
    .RX_CLKMUX_EN                       ( 1'b1),                                                
    .TX_XCLK_SEL                        ("TXUSR"),                                              
    .RX_XCLK_SEL                        ("RXDES"),   
    .TXOUT_DIV                          (OUT_DIV), 
    .RXOUT_DIV                          (OUT_DIV), 
    .LOCAL_MASTER                       (LOCAL_MASTER),   
    .RX_CLK_SLIP_OVRD                   ( 5'b00000),  
    .RXPMACLK_SEL                       ("DATA"),                                                                                                                           
    .USE_PCS_CLK_PHASE_SEL              ( 1'b0),           
   
    //----------------------------------------------------------------------------------------------     
    //  Programmable Divider Attributes
    //----------------------------------------------------------------------------------------------                                                                                                                       
    .TX_PROGCLK_SEL                     ("CPLL"),                               
    .TX_PROGDIV_CFG                     (PROGDIV_CFG),                      
    .RX_PROGDIV_CFG                     (PROGDIV_CFG),   
    .TX_PROGDIV_RATE                    (16'h0001),                          
    .RX_PROGDIV_RATE                    (16'h0001),                                   
               
    //----------------------------------------------------------------------------------------------
    //  CPLL Attributes
    //----------------------------------------------------------------------------------------------                 
    .CPLL_CFG0                          (16'h00FA), //(16'h20FA),               // Optimize for PCIe PLL compliance  
    .CPLL_CFG1                          (16'h0023), //(16'h24AA),          
    .CPLL_CFG2                          (16'h0002),                             
    .CPLL_CFG3                          ( 6'h00),  
    .CPLL_FBDIV                         (CPLL_FBDIV),  
    .CPLL_FBDIV_45                      (CPLL_FBDIV_45),    
    .CPLL_INIT_CFG0                     (16'h02B2),                
    .CPLL_LOCK_CFG                      (16'h01E8), //(16'h01E8),                             
    .CPLL_REFCLK_DIV                    ( 1),     
             
    //----------------------------------------------------------------------------------------------
    //  Reset Attributes
    //----------------------------------------------------------------------------------------------                
    .RESET_POWERSAVE_DISABLE            ( 1'b0),   
                                                                              
    //----------------------------------------------------------------------------------------------
    //  Reset Time Attributes
    //----------------------------------------------------------------------------------------------    
    .TX_DIVRESET_TIME                   ( 5'b00010), //( 5'b00001),  
    .TXPCSRESET_TIME	                  ( 5'b00011),
    .TXPMARESET_TIME	                  ( 5'b00011),
    .RX_DIVRESET_TIME                   ( 5'b00010), //( 5'b00001),  
    .RXBUFRESET_TIME                    ( 5'b00011),
    .RXCDRFREQRESET_TIME                ( 5'b10000), //( 5'b00001),  
    .RXCDRPHRESET_TIME                  ( 5'b00001),    
    .RXDFELPMRESET_TIME                 ( 7'b0001111),    
    .RXISCANRESET_TIME	                ( 5'b00001), 
    .RXOSCALRESET_TIME	                ( 5'b00011), 
    .RXPCSRESET_TIME	                  ( 5'b00011),   
    .RXPMARESET_TIME	                  ( 5'b00011),   
               
    //----------------------------------------------------------------------------------------------
    //  PCIe Attributes
    //----------------------------------------------------------------------------------------------
    .PCIE_BUFG_DIV_CTRL                 (PCIE_BUFG_DIV_CTRL),                  
    .PCIE_RXPCS_CFG_GEN3                (PCIE_RXPCS_CFG_GEN3),                 
    .PCIE_RXPMA_CFG                     (PCIE_PMA_CFG),                        
    .PCIE_TXPCS_CFG_GEN3                (PCIE_TXPCS_CFG_GEN3),                 
    .PCIE_TXPMA_CFG                     (PCIE_PMA_CFG),                        
    .PCS_PCIE_EN                        (PCS_PCIE_EN),  
    .PCIE_PLL_SEL_MODE_GEN12            (PCIE_PLL_SEL_MODE_GEN12),                  
    .PCIE_PLL_SEL_MODE_GEN3             (PCIE_PLL_SEL_MODE_GEN3),  
    .PCIE_PLL_SEL_MODE_GEN4             (PCIE_PLL_SEL_MODE_GEN4),                     
           
    //---------------------------------------------------------------------------------------------- 
    //  Data Width Attributes
    //----------------------------------------------------------------------------------------------                          
    .TX_DATA_WIDTH                      (20),                                                                                                                                         
    .RX_DATA_WIDTH                      (20),  
    .TX_INT_DATAWIDTH                   ( 0),                                                                
    .RX_INT_DATAWIDTH                   ( 0),   
    .TX_FABINT_USRCLK_FLOP              ( 1'b0), 
    .RX_FABINT_USRCLK_FLOP              ( 1'b0),                                                    
              
    //----------------------------------------------------------------------------------------------
    //  Analog Front End Attributes
    //----------------------------------------------------------------------------------------------
    .LPBK_BIAS_CTRL	                    ( 3'b100),                           
    .LPBK_EN_RCAL_B	                    ( 1'b0),                             
    .LPBK_EXT_RCAL	                    ( 4'b1000),                          
    .LPBK_RG_CTRL	                      ( 4'b1110),                             
    .RX_AFE_CM_EN                       ( 1'b0),
    .RX_BIAS_CFG0                       (16'h1554),
    .RX_CM_BUF_CFG                      ( 4'b1010),
    .RX_CM_BUF_PD                       ( 1'b0),                                           
    .RX_CM_SEL                          (RX_CM_SEL),                                                        
    .RX_CM_TRIM                         (10),    
    .RX_TUNE_AFE_OS                     ( 2'b00),
    .TERM_RCAL_CFG                      (15'b100001000010001),                                     
    .TERM_RCAL_OVRD                     ( 3'b000),             
                                                                                                    
    //----------------------------------------------------------------------------------------------  
    //  Receiver Detection Attributes
    //----------------------------------------------------------------------------------------------                                      
    .TX_RXDETECT_CFG                    (14'h0032),                                                      
    .TX_RXDETECT_REF                    (3),                                  
    
    //----------------------------------------------------------------------------------------------  
    //  TX Electrical Idle Attributes
    //----------------------------------------------------------------------------------------------   
    .TX_EIDLE_ASSERT_DELAY              (TX_EIDLE_ASSERT_DELAY),                            
    .TX_EIDLE_DEASSERT_DELAY            (TX_EIDLE_DEASSERT_DELAY),             
    .TX_IDLE_DATA_ZERO                  ( 1'b0),                                // Optimized for PCIe      
 
    //----------------------------------------------------------------------------------------------  
    //  RX OOB Attributes
    //----------------------------------------------------------------------------------------------   
    .OOB_PWRUP                          ( 1'b1),                                
    .OOBDIVCTL                          (OOBDIVCTL),                                            
    .RX_SIG_VALID_DLY                   ( 4),                                   // Optimized for PCIe
    .RXOOB_CFG                          ( 9'b000000110),                          
    .RXOOB_CLK_CFG                      ("PMA"),      
    
    //----------------------------------------------------------------------------------------------  
    //  RX Electrical Idle Attributes
    //----------------------------------------------------------------------------------------------                                                   
    .RX_DFE_LPM_HOLD_DURING_EIDLE       ( 1'b0),                                
    .RXBUF_EIDLE_HI_CNT                 ( 4'b0100),                             // Optimized for PCIe
    .RXBUF_EIDLE_LO_CNT                 ( 4'b0000),
    .RXBUF_RESET_ON_EIDLE               ("TRUE"),
    .RXCDR_FR_RESET_ON_EIDLE            ( 1'b0),
    .RXCDR_PH_RESET_ON_EIDLE            ( 1'b0),
    .RXCDR_HOLD_DURING_EIDLE            ( 1'b0),                                // Optimized for PCIe
    .RXELECIDLE_CFG                     ("SIGCFG_1"),                           // Optimized for PCIe
 
    //----------------------------------------------------------------------------------------------  
    //  Power Down Attributes
    //----------------------------------------------------------------------------------------------   
    .PD_TRANS_TIME_FROM_P2              (12'h03C),                                                     
    .PD_TRANS_TIME_NONE_P2              ( 8'h19),                                                      
    .PD_TRANS_TIME_TO_P2                ( 8'h64),   
    .TX_PMA_POWER_SAVE                  ( 1'b0),   
    .RX_PMA_POWER_SAVE                  ( 1'b0),                               
  
    //----------------------------------------------------------------------------------------------  
    //  Rate Change Attributes
    //---------------------------------------------------------------------------------------------- 
    .RATE_SW_USE_DRP                    ( 1'b0),                                // Advance PCIe feature
    .TRANS_TIME_RATE                    ( 8'h0E),             
    .TXBUF_RESET_ON_RATE_CHANGE         ("TRUE"),                              
    .RXBUF_RESET_ON_RATE_CHANGE         ("TRUE"),                              

    //----------------------------------------------------------------------------------------------
    //  TX Driver Attributes
    //----------------------------------------------------------------------------------------------                                   
    .TX_DEEMPH0                         ( 6'b010100),                           // -6.0 dB 
    .TX_DEEMPH1                         ( 6'b001101),                           // -3.5 dB
    .TX_DEEMPH2                         ( 6'b000000),                           //  0.0 dB 
    .TX_DEEMPH3                         ( 6'b000000),                           //  0.0 dB  
    .TX_DRIVE_MODE                      ("PIPE"),                                
    .TX_LOOPBACK_DRIVE_HIZ              ("FALSE"),                   
    .TX_MAINCURSOR_SEL                  ( 1'b0),   
    .TX_MARGIN_FULL_0                   ( 7'b1001111),                          // 1200 mV
    .TX_MARGIN_FULL_1                   ( 7'b1001110),                          // 1100 mV
    .TX_MARGIN_FULL_2                   ( 7'b1001100),                          // 1000 mV 
    .TX_MARGIN_FULL_3                   ( 7'b1001010),                          //  900 mV
    .TX_MARGIN_FULL_4                   ( 7'b1001000),                          //  800 mV
    .TX_MARGIN_LOW_0                    ( 7'b1000110),                          //  700 mV            
    .TX_MARGIN_LOW_1                    ( 7'b1000101),                          //  600 mV           
    .TX_MARGIN_LOW_2                    ( 7'b1000011),                          //  500 mV          
    .TX_MARGIN_LOW_3                    ( 7'b1000010),                          //  400 mV           
    .TX_MARGIN_LOW_4                    ( 7'b1000000),                          //  300 mV                               
   
    //----------------------------------------------------------------------------------------------    
    //  Comma Align & Detect Attributes
    //----------------------------------------------------------------------------------------------       
    .ALIGN_COMMA_DOUBLE                 (ALIGN_COMMA_DOUBLE),                                                  
    .ALIGN_COMMA_ENABLE                 (10'b1111111111),                                           
    .ALIGN_COMMA_WORD                   ( 1),                                                       
    .ALIGN_MCOMMA_DET                   ("TRUE"),                                                   
    .ALIGN_MCOMMA_VALUE                 (10'b1010000011),                                           
    .ALIGN_PCOMMA_DET                   ("TRUE"),                                                   
    .ALIGN_PCOMMA_VALUE                 (10'b0101111100),                                           
    .DEC_MCOMMA_DETECT                  ("TRUE"),                                                      
    .DEC_PCOMMA_DETECT                  ("TRUE"),                                                      
    .DEC_VALID_COMMA_ONLY               ("FALSE"),                                                     
    .SHOW_REALIGN_COMMA                 (SHOW_REALIGN_COMMA),       
   
    //----------------------------------------------------------------------------------------------   
    //  8B/10B Attributes                                                                             
    //----------------------------------------------------------------------------------------------                   
    .RX_DISPERR_SEQ_MATCH               ("TRUE"),        
   
    //----------------------------------------------------------------------------------------------  
    //  TX Buffer Attributes
    //----------------------------------------------------------------------------------------------                      
    .TX_FIFO_BYP_EN                     ( 1'b1),                                
    .TXBUF_EN                           ("FALSE"),        
    .TXFIFO_ADDR_CFG                    ("LOW"),                                                                                      
 
    //----------------------------------------------------------------------------------------------
    //  RX Buffer Attributes                                                                        
    //----------------------------------------------------------------------------------------------     
    .RXBUF_ADDR_MODE                    ("FULL"),                               
    .RXBUF_EN                           ("TRUE"),
    .RXBUF_RESET_ON_CB_CHANGE           ("TRUE"),
    .RXBUF_RESET_ON_COMMAALIGN          ("FALSE"),
    .RXBUF_THRESH_OVFLW                 (RXBUF_THRESH_OVFLW),                                                      
    .RXBUF_THRESH_OVRD                  ("TRUE"),                             
    .RXBUF_THRESH_UNDFLW                (RXBUF_THRESH_UNDFLW),                                    
    .RX_BUFFER_CFG                      ( 6'b000000),
    .RX_DEFER_RESET_BUF_EN              ("TRUE"), 
   
    //----------------------------------------------------------------------------------------------   
    //  PCIe Gen3 RX Buffer Attributes                                                                                   
    //----------------------------------------------------------------------------------------------   
    .PCI3_AUTO_REALIGN                  ("OVR_1K_BLK"),                           
    .PCI3_PIPE_RX_ELECIDLE              ( 1'b0),                                
    .PCI3_RX_ASYNC_EBUF_BYPASS          ( 2'b00),                               
    .PCI3_RX_ELECIDLE_EI2_ENABLE        ( 1'b0),                                
    .PCI3_RX_ELECIDLE_H2L_COUNT         ( 6'b000000),                           
    .PCI3_RX_ELECIDLE_H2L_DISABLE       ( 3'b000),                              
    .PCI3_RX_ELECIDLE_HI_COUNT          ( 6'b000000),                           
    .PCI3_RX_ELECIDLE_LP4_DISABLE       ( 1'b0),                                
    .PCI3_RX_FIFO_DISABLE               ( 1'b0),                                
       
    //----------------------------------------------------------------------------------------------   
    //  PCIe Gen3 Clock Correction Attributes                                                                                   
    //----------------------------------------------------------------------------------------------          
    .PCIE3_CLK_COR_EMPTY_THRSH          (PCIE3_CLK_COR_EMPTY_THRSH),                           
    .PCIE3_CLK_COR_FULL_THRSH           (PCIE3_CLK_COR_FULL_THRSH),                          
    .PCIE3_CLK_COR_MAX_LAT              (PCIE3_CLK_COR_MAX_LAT),                          
    .PCIE3_CLK_COR_MIN_LAT              (PCIE3_CLK_COR_MIN_LAT),                          
    .PCIE3_CLK_COR_THRSH_TIMER          (PCIE3_CLK_COR_THRSH_TIMER),                      
       
    //---------------------------------------------------------------------------------------------- 
    //  Clock Correction Attributes
    //----------------------------------------------------------------------------------------------             
    .CBCC_DATA_SOURCE_SEL               ("DECODED"),  
    .CLK_COR_KEEP_IDLE                  (CLK_COR_KEEP_IDLE),
    .CLK_COR_MAX_LAT                    (CLK_COR_MAX_LAT),                                   
    .CLK_COR_MIN_LAT                    (CLK_COR_MIN_LAT),                                  
    .CLK_COR_PRECEDENCE                 ("TRUE"),
    .CLK_COR_REPEAT_WAIT                (0),
    .CLK_COR_SEQ_1_1                    (CLK_COR_SEQ_1_1),
    .CLK_COR_SEQ_1_2                    (CLK_COR_SEQ_1_2),
    .CLK_COR_SEQ_1_3                    (10'b0000000000),
    .CLK_COR_SEQ_1_4                    (10'b0000000000),
    .CLK_COR_SEQ_1_ENABLE               (4'b1111),
    .CLK_COR_SEQ_2_1                    (10'b0000000000),
    .CLK_COR_SEQ_2_2                    (10'b0000000000),
    .CLK_COR_SEQ_2_3                    (10'b0000000000),
    .CLK_COR_SEQ_2_4                    (10'b0000000000),
    .CLK_COR_SEQ_2_ENABLE               (CLK_COR_SEQ_2_ENABLE),
    .CLK_COR_SEQ_2_USE                  ("FALSE"),
    .CLK_COR_SEQ_LEN                    (CLK_COR_SEQ_LEN),
    .CLK_CORRECT_USE                    ("TRUE"),                
       
    //---------------------------------------------------------------------------------------------- 
    //  FTS Deskew Attributes                                                                            
    //----------------------------------------------------------------------------------------------                                         
    .FTS_DESKEW_SEQ_ENABLE              ( 4'b1111),                                        
    .FTS_LANE_DESKEW_CFG                ( 4'b1111),                                          
    .FTS_LANE_DESKEW_EN                 ("FALSE"),           
       
    //---------------------------------------------------------------------------------------------- 
    //  Channel Bonding Attributes (Disabled)
    //----------------------------------------------------------------------------------------------          
    .CHAN_BOND_KEEP_ALIGN               ("FALSE"),
    .CHAN_BOND_MAX_SKEW                 ( 1),
    .CHAN_BOND_SEQ_1_1                  (10'b0000000000),
    .CHAN_BOND_SEQ_1_2                  (10'b0000000000),
    .CHAN_BOND_SEQ_1_3                  (10'b0000000000),
    .CHAN_BOND_SEQ_1_4                  (10'b0000000000),
    .CHAN_BOND_SEQ_1_ENABLE             ( 4'b1111),
    .CHAN_BOND_SEQ_2_1                  (10'b0000000000),
    .CHAN_BOND_SEQ_2_2                  (10'b0000000000),
    .CHAN_BOND_SEQ_2_3                  (10'b0000000000),
    .CHAN_BOND_SEQ_2_4                  (10'b0000000000),  
    .CHAN_BOND_SEQ_2_ENABLE             ( 4'b1111),
    .CHAN_BOND_SEQ_2_USE                ("FALSE"), 
    .CHAN_BOND_SEQ_LEN                  ( 1),                                                           
  
    //----------------------------------------------------------------------------------------------            
    //  TX Sync Alignment Attributes                                                                              
    //----------------------------------------------------------------------------------------------     
    .TXDLY_CFG                          (16'b1000000000010000),    
    .TXDLY_LCFG                         (16'b0000000000110000),                
    .TXPH_CFG                           (16'b0000000100100011), //(16'b0000000100000011),               
    .TXPH_CFG2                          (16'b0000000000000000),                 
    .TXPH_MONITOR_SEL                   ( 5'b00000),
    .TXPHDLY_CFG0                       (16'b0110000000100000),                 
    .TXPHDLY_CFG1                       (16'b0000000000000010),              
                                                                                    
    //----------------------------------------------------------------------------------------------            
    //  TX Auto Sync Alignment Attributes                                                                               
    //----------------------------------------------------------------------------------------------                
    .TXSYNC_MULTILANE                   (MULTI_LANE),                                                                                                              
    .TXSYNC_OVRD                        (1'b0),                                 // Select auto TXSYNC mode                                                                                 
    .TXSYNC_SKIP_DA                     (1'b0),                     
                                                                                                    
    //----------------------------------------------------------------------------------------------            
    //  RX Sync Alignment Attributes (Not used)                                                                             
    //----------------------------------------------------------------------------------------------    
  //.RXDLY_CFG                          (16'h001F),   
  //.RXDLY_LCFG                         (16'h0030),   
  //.RXPH_MONITOR_SEL                   (5'b00000),
  //.RXPHBEACON_CFG                     (16'h0000),
  //.RXPHDLY_CFG                        (16'h2020),
  //.RXPHSAMP_CFG                       (16'h2100),
  //.RXPHSLIP_CFG                       (16'h9933),                             
     
    //----------------------------------------------------------------------------------------------            
    //  RX Auto Sync Alignment Attributes (Not used)                                                                                
    //----------------------------------------------------------------------------------------------                
  //.RXSYNC_MULTILANE                   (1'b0),                                                                                                              
  //.RXSYNC_OVRD                        (1'b0),                                                                                         
  //.RXSYNC_SKIP_DA                     (1'b0),                   
  
    //----------------------------------------------------------------------------------------------  
    //  Gearbox Attributes (Not used)                                                                
    //---------------------------------------------------------------------------------------------- 
  //.GEARBOX_MODE                       ( 5'b00000), 
  //.TX_SAMPLE_PERIOD                   ( 3'b101),
  //.RX_SAMPLE_PERIOD                   ( 3'b101),
  //.TXGEARBOX_EN                       ("FALSE"),
  //.RXGEARBOX_EN                       ("FALSE"),    
  //.TXGBOX_FIFO_INIT_RD_ADDR           ( 4),
  //.RXGBOX_FIFO_INIT_RD_ADDR           ( 4),
  //.RXSLIDE_AUTO_WAIT                  ( 7),                                                         
    .RXSLIDE_MODE                       (RXSLIDE_MODE),                          

    //----------------------------------------------------------------------------------------------
    //  PCS Reserved Attributes
    //----------------------------------------------------------------------------------------------
    .PCS_RSVD0                          (PCS_RSVD0),
  
    //----------------------------------------------------------------------------------------------  
    //  PMA Reserved Attributes
    //----------------------------------------------------------------------------------------------      
    .TX_PMA_RSV0                        (16'b0000000000001000),                             
    .RX_PMA_RSV0                        (16'b0000000000000000),                                        
      
    //----------------------------------------------------------------------------------------------
    //  CFOK Attributes                                                                 
    //----------------------------------------------------------------------------------------------              
    .RXCFOK_CFG0                        (16'b0000000000000000), //(16'b0011111000000000),   
    .RXCFOK_CFG1                        (16'b1000000000010101), //(16'b0000000001000010),    
    .RXCFOK_CFG2                        (16'b0000001010101110), //(16'b0000000000101101),  

    //----------------------------------------------------------------------------------------------
    //  RX CTLE
    //----------------------------------------------------------------------------------------------  
    .CTLE3_OCAP_EXT_CTRL	              ( 3'b000),                           
    .CTLE3_OCAP_EXT_EN	                ( 1'b0),                                
    .RX_EN_CTLE_RCAL_B                  ( 1'b0),                              

    //----------------------------------------------------------------------------------------------    
    //  RX LPM Attributes
    //----------------------------------------------------------------------------------------------        
    .RXLPM_CFG                          (16'b0000_0000_0000_0000),    
    .RXLPM_GC_CFG                       (16'b1000_0000_0000_0000),
    .RXLPM_KH_CFG0                      (16'b0000_0000_0000_0000), //(16'b0000000000000000),    
    .RXLPM_KH_CFG1                      (16'b0000_0000_0000_0010), //(16'b0000000000000010),    
    .RXLPM_OS_CFG0                      (16'b0000_0000_0000_0000),
    .RXLPM_OS_CFG1                      (16'b1000_0000_0000_0010), //(16'b0000000000000000), 
 
    //----------------------------------------------------------------------------------------------    
    //  RX DFE Attributes
    //----------------------------------------------------------------------------------------------       
    .RXDFE_CFG0                         (16'b0000101000000000), //(16'b0000110000000000),    
    .RXDFE_CFG1                         (16'b0000001010000000),
    .RXDFE_GC_CFG0                      (16'b0000000000000000), //(16'b0001111000000000),    
    .RXDFE_GC_CFG1                      (16'b1000000000000000), //(16'h1900),   different from GTY             
    .RXDFE_GC_CFG2                      (16'b1111111111100000), //(16'h0000),   different from GTY             
    .RXDFE_H2_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_H2_CFG1                      (16'b0000000000000010), //(16'b0000000000000010),    
    .RXDFE_H3_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_H3_CFG1                      (16'b1000000000000010), //(16'b0000000000000010),    
    .RXDFE_H4_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_H4_CFG1                      (16'b1000000000000010), //(16'b0000000000000011),    
    .RXDFE_H5_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_H5_CFG1                      (16'b1000000000000010), //(16'b0000000000000010),    
    .RXDFE_H6_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_H6_CFG1                      (16'b1000000000000010), //(16'b0000000000000010),    
    .RXDFE_H7_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_H7_CFG1                      (16'b1000000000000010), //(16'b0000000000000010),    
    .RXDFE_H8_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_H8_CFG1                      (16'b1000000000000010), //(16'b0000000000000010),    
    .RXDFE_H9_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_H9_CFG1                      (16'b1000000000000010), //(16'b0000000000000010),    
    .RXDFE_HA_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_HA_CFG1                      (16'b1000000000000010), //(16'b0000000000000010),    
    .RXDFE_HB_CFG0                      (16'b0000000000000000), //(16'b0010000000000000),    
    .RXDFE_HB_CFG1                      (16'b1000000000000010), //(16'b0000000000000010),    
    .RXDFE_HC_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_HC_CFG1                      (16'b1000000000000010), //(16'b0000000000000010),    
    .RXDFE_HD_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_HD_CFG1                      (16'b1000000000000010), //(16'b0000000000000010),    
    .RXDFE_HE_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_HE_CFG1                      (16'b1000000000000010), //(16'b0000000000000010),    
    .RXDFE_HF_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_HF_CFG1                      (16'b1000000000000010), //(16'b0000000000000010),    
    .RXDFE_OS_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_OS_CFG1                      (16'b1000000000000010), //(16'b0000001000000000),    
    .RXDFE_PWR_SAVING                   (RXDFE_PWR_SAVING),
    .RXDFE_UT_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_UT_CFG1                      (16'b0000000000000011), //(16'b0000000000000010),    
    .RXDFE_UT_CFG2                      (16'b0000000000000000),
    .RXDFE_VP_CFG0                      (16'b0000000000000000), //(16'b0000000000000000),    
    .RXDFE_VP_CFG1                      (16'b1000000000110011), //(16'b0000000000100010),    
    .RXDFELPM_KL_CFG0                   (16'b0000000000000000),                  
    .RXDFELPM_KL_CFG1                   (16'b1010000011100010),             
    .RXDFELPM_KL_CFG2                   (16'b0000000100000000),                        
    .RX_DFE_AGC_CFG0                    ( 2'b10),                               
    .RX_DFE_AGC_CFG1                    ( 4),  
    .RX_DFE_KL_LPM_KH_CFG0              ( 1),
    .RX_DFE_KL_LPM_KH_CFG1              ( 4),
    .RX_DFE_KL_LPM_KL_CFG0              ( 2'b01),
    .RX_DFE_KL_LPM_KL_CFG1              ( 4),   
    .RX_DFELPM_CFG0                     ( 6),                                                            
    .RX_DFELPM_CFG1                     ( 1'b1),                                                               
    .RX_DFELPM_KLKH_AGC_STUP_EN         ( 1'b1),   
          
    //----------------------------------------------------------------------------------------------  
    //  TX PI attributes
    //----------------------------------------------------------------------------------------------
    .TX_PHICAL_CFG0	                    (16'h0000),                           
    .TX_PHICAL_CFG1	                    (16'h7e00),
    .TX_PHICAL_CFG2	                    (16'h0200), //(16'h0000),  
    .TX_PI_BIASSET	                    (TX_PI_BIASSET),                                  
    .TXPI_CFG0                          ( 2'b00),
    .TXPI_CFG1                          ( 2'b00),
    .TXPI_CFG2                          ( 2'b00),
    .TXPI_CFG3                          ( 1'b0),
    .TXPI_CFG4                          ( 1'b0),
    .TXPI_CFG5                          ( 3'b000),
    .TXPI_GRAY_SEL                      ( 1'b0),
    .TXPI_INVSTROBE_SEL                 ( 1'b0),
    .TXPI_LPM                           ( 1'b0),
    .TXPI_PPM_CFG                       ( 8'b00000000),
    .TXPI_PPMCLK_SEL                    ("TXUSRCLK2"),
    .TXPI_SYNFREQ_PPM                   ( 3'b001),
    .TXPI_VREFSEL                       ( 1'b0),
    
    //----------------------------------------------------------------------------------------------  
    //  RX PI Attributes
    //----------------------------------------------------------------------------------------------    
    .RXPI_AUTO_BW_SEL_BYPASS            ( 1'b0),
    .RXPI_CFG0                          (RXPI_CFG0),
    .RXPI_CFG1                          (16'h0000),
    .RXPI_LPM                           ( 1'b0),
    .RXPI_SEL_LC                        ( 2'b00),
    .RXPI_STARTCODE                     ( 2'b00),
    .RXPI_VREFSEL                       ( 1'b0),              

    //----------------------------------------------------------------------------------------------
    //  RX CDR Attributes
    //----------------------------------------------------------------------------------------------    
    .CDR_SWAP_MODE_EN                   ( 1'b0),                 
    .RX_WIDEMODE_CDR                    ( 2'b00),                               //Gen1/2 wide mode    
    .RX_WIDEMODE_CDR_GEN3               ( 2'b00), 
    .RX_WIDEMODE_CDR_GEN4               ( 2'b01),
    .RXCDR_CFG0                         (RXCDR_CFG0), 
    .RXCDR_CFG0_GEN3                    (RXCDR_CFG0_GEN3), 
    .RXCDR_CFG1                         (RXCDR_CFG1), 
    .RXCDR_CFG1_GEN3                    (RXCDR_CFG1_GEN3), 
    .RXCDR_CFG2                         (RXCDR_CFG2), 
    .RXCDR_CFG2_GEN3                    (RXCDR_CFG2_GEN3), 
    .RXCDR_CFG2_GEN4                    (RXCDR_CFG2_GEN4), 
    .RXCDR_CFG3                         (RXCDR_CFG3), 
    .RXCDR_CFG3_GEN3                    (RXCDR_CFG3_GEN3), 
    .RXCDR_CFG3_GEN4                    (RXCDR_CFG3_GEN4),
    .RXCDR_CFG4                         (RXCDR_CFG4), 
    .RXCDR_CFG4_GEN3                    (RXCDR_CFG4_GEN3), 
    .RXCDR_CFG5                         (RXCDR_CFG5), 
    .RXCDR_CFG5_GEN3                    (RXCDR_CFG5_GEN3), 
    .RXCDR_LOCK_CFG0                    (16'b0001_0010_0000_0001), //(16'h0001),  
    .RXCDR_LOCK_CFG1                    (16'b1001_1111_1111_1111), //(16'h0000),  
    .RXCDR_LOCK_CFG2                    (16'b0111_0111_1100_0011), //(16'b0000),  
    .RXCDR_LOCK_CFG3                    (16'b0000_0000_0000_0001), //(16'h0000),  

    //---------------------------------------------------------------------------------------------- 
    //  Eye Scan Attributes
    //----------------------------------------------------------------------------------------------
    .ES_CLK_PHASE_SEL                   ( 1'b0),                           
    .ES_CONTROL                         ( 6'b000000),                      
    .ES_ERRDET_EN                       ("FALSE"),                        
    .ES_EYE_SCAN_EN                     ("FALSE"),                        
    .ES_HORZ_OFFSET                     (12'b000000000000),                       
    .ES_PRESCALE                        ( 5'b00000),                                
    .ES_QUAL_MASK0                      (16'b0000000000000000),           
    .ES_QUAL_MASK1                      (16'b0000000000000000),           
    .ES_QUAL_MASK2                      (16'b0000000000000000),           
    .ES_QUAL_MASK3                      (16'b0000000000000000),           
    .ES_QUAL_MASK4                      (16'b0000000000000000),       
    .ES_QUAL_MASK5                      (16'b0000000000000000),           
    .ES_QUAL_MASK6                      (16'b0000000000000000),           
    .ES_QUAL_MASK7                      (16'b0000000000000000),           
    .ES_QUAL_MASK8                      (16'b0000000000000000),           
    .ES_QUAL_MASK9                      (16'b0000000000000000),         
    .ES_QUALIFIER0                      (16'b0000000000000000),           
    .ES_QUALIFIER1                      (16'b0000000000000000),           
    .ES_QUALIFIER2                      (16'b0000000000000000),           
    .ES_QUALIFIER3                      (16'b0000000000000000),           
    .ES_QUALIFIER4                      (16'b0000000000000000), 
    .ES_QUALIFIER5                      (16'b0000000000000000),           
    .ES_QUALIFIER6                      (16'b0000000000000000),           
    .ES_QUALIFIER7                      (16'b0000000000000000),           
    .ES_QUALIFIER8                      (16'b0000000000000000),           
    .ES_QUALIFIER9                      (16'b0000000000000000),   
    .ES_SDATA_MASK0                     (16'b0000000000000000),           
    .ES_SDATA_MASK1                     (16'b0000000000000000),           
    .ES_SDATA_MASK2                     (16'b0000000000000000),           
    .ES_SDATA_MASK3                     (16'b0000000000000000),           
    .ES_SDATA_MASK4                     (16'b0000000000000000), 
    .ES_SDATA_MASK5                     (16'b0000000000000000),           
    .ES_SDATA_MASK6                     (16'b0000000000000000),           
    .ES_SDATA_MASK7                     (16'b0000000000000000),           
    .ES_SDATA_MASK8                     (16'b0000000000000000),   
    .ES_SDATA_MASK9                     (16'b0000000000000000),          
    .EYE_SCAN_SWAP_EN                   ( 1'b0),
    .RX_EYESCAN_VS_CODE                 ( 7'b0000000),
    .RX_EYESCAN_VS_NEG_DIR              ( 1'b0),
    .RX_EYESCAN_VS_RANGE                ( 2'b00),
    .RX_EYESCAN_VS_UT_SIGN              ( 1'b0),                        
  
    //----------------------------------------------------------------------------------------------
    //  Loopback & PRBS Attributes
    //----------------------------------------------------------------------------------------------
    .RXPRBS_ERR_LOOPBACK                ( 1'b0),     
    .RXPRBS_LINKACQ_CNT                 (15),                                                   

    //----------------------------------------------------------------------------------------------   
    //  Digital Monitor Attribute
    //----------------------------------------------------------------------------------------------                     
    .DMONITOR_CFG0                      (10'b0000000000),                                                  
    .DMONITOR_CFG1                      ( 8'b00000000),                                                   

    //----------------------------------------------------------------------------------------------   
    //  AC JTAG Attributes
    //----------------------------------------------------------------------------------------------                     
    .ACJTAG_DEBUG_MODE                  ( 1'b0),                                                        
    .ACJTAG_MODE                        ( 1'b0),                                                        
    .ACJTAG_RESET                       ( 1'b0),      
    
    //----------------------------------------------------------------------------------------------
    //  USB Attributes
    //----------------------------------------------------------------------------------------------                 
    .USB_BOTH_BURST_IDLE                ( 1'b0),
    .USB_BURSTMAX_U3WAKE	              ( 7'b1111111),
    .USB_BURSTMIN_U3WAKE	              ( 7'b1100011),
    .USB_CLK_COR_EQ_EN                  ( 1'b1),                              
    .USB_EXT_CNTL                       ( 1'b1),
    .USB_IDLEMAX_POLLING                (10'b1010111011),
    .USB_IDLEMIN_POLLING                (10'b0100101011),
    .USB_LFPS_TPERIOD	                  ( 4'b0011),
    .USB_LFPS_TPERIOD_ACCURATE	        ( 1'b1),
    .USB_LFPSPING_BURST	                ( 9'b000000101),
    .USB_LFPSPOLLING_BURST	            ( 9'b000110001),
    .USB_LFPSPOLLING_IDLE_MS	          ( 9'b000000100),
    .USB_LFPSU1EXIT_BURST	              ( 9'b000011101),
    .USB_LFPSU2LPEXIT_BURST_MS	        ( 9'b001100011),
    .USB_LFPSU3WAKE_BURST_MS	          ( 9'b111110011),
    .USB_MODE                           (USB_MODE), 
    .USB_PCIE_ERR_REP_DIS               ( 1'b0),                                // For PCIe Debug
    .USB_PING_SATA_MAX_INIT             (21),
    .USB_PING_SATA_MIN_INIT             (12),
    .USB_POLL_SATA_MAX_BURST            ( 8),
    .USB_POLL_SATA_MIN_BURST            ( 4),
    .USB_RAW_ELEC                       ( 1'b1),                               
    .USB_RXIDLE_P0_CTRL                 ( 1'b1),
    .USB_TXIDLE_TUNE_ENABLE             ( 1'b1),
    .USB_U1_SATA_MAX_WAKE               ( 7),
    .USB_U1_SATA_MIN_WAKE               ( 4),
    .USB_U2_SAS_MAX_COM                 (64),   
    .USB_U2_SAS_MIN_COM                 (36),
    
    //---------------------------------------------------------------------------------------------- 
    //  SAS & SATA Attributes (Not used)
    //---------------------------------------------------------------------------------------------- 
  //.SAS12G_MODE                        ( 1'b0),
  //.SATA_BURST_SEQ_LEN                 ( 4'b1111),
  //.SATA_BURST_VAL                     ( 3'b100),
  //.SATA_CPLL_CFG                      ("VCO_3000MHZ"),
  //.SATA_EIDLE_VAL                     ( 3'b100), 
            
    //---------------------------------------------------------------------------------------------- 
    //  CKCAL Attributes
    //---------------------------------------------------------------------------------------------- 
    .CKCAL1_CFG_0	                      (16'hC0C0), //(16'b0000000000000000), 
    .CKCAL1_CFG_1	                      (16'h50C0), //(16'b0000000000000000), 
    .CKCAL1_CFG_2	                      (16'b0000000000001010),
    .CKCAL1_CFG_3	                      (16'b0000000000000000),
    .CKCAL2_CFG_0	                      (16'hC0C0), //(16'b0000000000000000), 
    .CKCAL2_CFG_1	                      (16'h80C0), //(16'b0000000000000000), 
    .CKCAL2_CFG_2	                      (16'b0000000000000000),
    .CKCAL2_CFG_3	                      (16'b0000000000000000),
    .CKCAL2_CFG_4	                      (16'b0000000000000000),
    .CKCAL_RSVD0	                      (16'h0000),
    .CKCAL_RSVD1	                      (16'b0000010000000000), //(16'h0000),
    .RXCKCAL1_I_LOOP_RST_CFG	          (16'h0004),
    .RXCKCAL1_IQ_LOOP_RST_CFG	          (16'h0004),
    .RXCKCAL1_Q_LOOP_RST_CFG	          (16'h0004),
    .RXCKCAL2_D_LOOP_RST_CFG	          (16'h0004),
    .RXCKCAL2_DX_LOOP_RST_CFG	          (16'h0004),
    .RXCKCAL2_S_LOOP_RST_CFG	          (16'h0004),
    .RXCKCAL2_X_LOOP_RST_CFG	          (16'h0004),
  
    //----------------------------------------------------------------------------------------------
    //  Summer Attributes
    //----------------------------------------------------------------------------------------------
    .RX_SUM_DFETAPREP_EN                ( 1'b0),
    .RX_SUM_IREF_TUNE                   (RX_SUM_IREF_TUNE),
    .RX_SUM_VCM_OVWR                    ( 1'b0),
    .RX_SUM_VCMTUNE                     (RX_SUM_VCMTUNE),
    .RX_SUM_VREF_TUNE                   ( 3'b100),

    //----------------------------------------------------------------------------------------------
    //  Attributes
    //----------------------------------------------------------------------------------------------                 
    .A_RXOSCALRESET                     ( 1'b0),   
    .A_RXPROGDIVRESET                   ( 1'b0),
    .A_RXTERMINATION                    ( 1'b1),
    .A_TXDIFFCTRL                       ( 5'b11111),
    .A_TXPROGDIVRESET                   ( 1'b0),
    .ADAPT_CFG0                         (16'b0001000000000000), //(16'b1001001000000000),   
    .ADAPT_CFG1                         (16'b1100101100000000), //(16'b1000000000011100),   
    .ADAPT_CFG2                         (16'b0000000000000000),   
    .CAPBYPASS_FORCE                    ( 1'b0),                                
    .CH_HSPMUX                          (16'b0110_1101_0110_1101), //(16'h0000),   
    .DDI_CTRL                           ( 2'b00),
    .DDI_REALIGN_WAIT                   (15),
    .DELAY_ELEC                         ( 1'b0),                                
    .ISCAN_CK_PH_SEL2                   ( 1'b0),                                
    .PREIQ_FREQ_BST                     ( 1),                                   
    .PROCESS_PAR                        ( 3'b010), 
    .RX_CAPFF_SARC_ENB                  ( 1'b0),    
    .RX_DDI_SEL                         ( 6'b000000),  
    .RX_DEGEN_CTRL                      ( 3'b011),                              
    .RX_DIV2_MODE_B                     ( 1'b0),                                
    .RX_EN_HI_LR                        ( 1'b1),
    .RX_EXT_RL_CTRL                     ( 9'b000000000),                        
    .RX_RESLOAD_CTRL	                  ( 4'b0000),                             
    .RX_RESLOAD_OVRD	                  ( 1'b0),                                
    .RX_VREG_CTRL	                      ( 3'b101),                              
    .RX_VREG_PDB	                      ( 1'b1),                                
    .RX_XMODE_SEL	                      ( 1'b0),                                
    .TAPDLY_SET_TX                      ( 2'b00),
    .TEMPERATURE_PAR                    ( 4'b0010),
    .TST_RSV0                           ( 8'b00000000),                                     
    .TST_RSV1                           ( 8'b00000000),
    .TX_DCC_LOOP_RST_CFG                (16'h0004),                             
    .TX_DRVMUX_CTRL                     ( 2),                                   
    .TX_PREDRV_CTRL                     ( 2),                                   
    .TX_PMADATA_OPT                     ( 1'b0)    
)                                                                                                   
gthe4_channel_smsw_i                                                                                     
(                                                                                                                                                                                                   
    //----------------------------------------------------------------------------------------------
    //  Clock Ports
    //----------------------------------------------------------------------------------------------
    .GTGREFCLK                          ( 1'd0),                                                     
    .GTREFCLK0                          (GT_GTREFCLK0),                                            
    .GTREFCLK1                          ( 1'd0),                                                    
    .GTNORTHREFCLK0                     ( 1'd0),                                                    
    .GTNORTHREFCLK1                     ( 1'd0),                                                    
    .GTSOUTHREFCLK0                     ( 1'd0),                                                    
    .GTSOUTHREFCLK1                     ( 1'd0),                                             
    .TXUSRCLK                           (GT_TXUSRCLK),                                              
    .RXUSRCLK                           (GT_RXUSRCLK),                                              
    .TXUSRCLK2                          (GT_TXUSRCLK2),                                             
    .RXUSRCLK2                          (GT_RXUSRCLK2),  
    .TXPLLCLKSEL                        (PLLCLKSEL),            
    .RXPLLCLKSEL                        (PLLCLKSEL),                                                    
    .TXSYSCLKSEL                        (SYSCLKSEL),                                             
    .RXSYSCLKSEL                        (SYSCLKSEL),                             
    .TXOUTCLKSEL                        (GT_TXOUTCLKSEL),                                // Select TXPROGDIVCLK
    .RXOUTCLKSEL                        ( 3'd2),                                // Select RXOUTCLKPMA
    .CLKRSVD0                           ( 1'd0),          
    .CLKRSVD1                           ( 1'd0),            
                                                                                                   
    .TXOUTCLK                           (GT_TXOUTCLK),                                             
    .RXOUTCLK                           (GT_RXOUTCLK),                                                        
    .TXOUTCLKFABRIC                     (GT_TXOUTCLKFABRIC),                                                        
    .RXOUTCLKFABRIC                     (GT_RXOUTCLKFABRIC),                                                        
    .TXOUTCLKPCS                        (GT_TXOUTCLKPCS),                                                        
    .RXOUTCLKPCS                        (GT_RXOUTCLKPCS),  
    .RXRECCLKOUT                        (GT_RXRECCLKOUT),                                                    
    .GTREFCLKMONITOR                    (),                                 
    
    //----------------------------------------------------------------------------------------------
    //  BUFG_GT Controller Ports
    //----------------------------------------------------------------------------------------------
    .BUFGTCE                            (GT_BUFGTCE),      
    .BUFGTCEMASK                        (GT_BUFGTCEMASK), 
    .BUFGTDIV                           (GT_BUFGTDIV), 
    .BUFGTRESET                         (GT_BUFGTRESET), 
    .BUFGTRSTMASK                       (GT_BUFGTRSTMASK),       
    
    //----------------------------------------------------------------------------------------------
    //  CPLL Ports
    //----------------------------------------------------------------------------------------------
    .CPLLFREQLOCK                       (GT_MASTER_CPLLLOCK),                 
    .CPLLLOCKDETCLK                     ( 1'd0),                              
    .CPLLLOCKEN                         ( 1'd1),    
    .CPLLPD                             (GT_CPLLPD),    
    .CPLLREFCLKSEL                      ( 3'd1),                               
    .CPLLRESET                          (GT_CPLLRESET),                               
  
    .CPLLFBCLKLOST                      (),     
    .CPLLLOCK                           (GT_CPLLLOCK),                                            
    .CPLLREFCLKLOST                     (),                    
             
    //----------------------------------------------------------------------------------------------
    //  QPLL Ports                                                                                   
    //----------------------------------------------------------------------------------------------
    .QPLL0CLK                           (GT_QPLL0CLK),                           
    .QPLL0REFCLK                        (GT_QPLL0REFCLK),                        
    .QPLL0FREQLOCK                      (GT_QPLL0LOCK),                         
    .QPLL1CLK                           (GT_QPLL1CLK),  
    .QPLL1REFCLK                        (GT_QPLL1REFCLK),           
    .QPLL1FREQLOCK                      (GT_QPLL1LOCK),                         
    
    //----------------------------------------------------------------------------------------------
    //  Reset Ports
    //----------------------------------------------------------------------------------------------                                                                                                                             
    .GTTXRESET                          (GT_GTTXRESET),                                             
    .GTRXRESET                          (GT_GTRXRESET),  
    .GTRXRESETSEL                       ( 1'd0),                                
    .GTTXRESETSEL                       ( 1'd0),                                
    .TXPROGDIVRESET                     (GT_TXPROGDIVRESET),                       
    .RXPROGDIVRESET                     ( 1'd0),                                                                            
    .TXPMARESET                         (GT_TXPMARESET),                                            
    .RXPMARESET                         (GT_RXPMARESET),                                            
    .TXPCSRESET                         (GT_TXPCSRESET),   
    .RXPCSRESET                         (GT_RXPCSRESET),   
    .TXUSERRDY                          (GT_TXUSERRDY),                                             
    .RXUSERRDY                          (GT_RXUSERRDY),   
    .CFGRESET                           ( 1'd0),                                                    
    .RESETOVRD                          (GT_RESETOVRD),  
    .RXOOBRESET                         ( 1'd0),                                              
                                           
    .GTPOWERGOOD                        (GT_GTPOWERGOOD), 
    .TXPRGDIVRESETDONE                  (GT_TXPROGDIVRESETDONE),
    .RXPRGDIVRESETDONE                  (),        
    .TXPMARESETDONE                     (GT_TXPMARESETDONE),    
    .RXPMARESETDONE                     (GT_RXPMARESETDONE),                                                                                                      
    .TXRESETDONE                        (GT_TXRESETDONE),                                           
    .RXRESETDONE                        (GT_RXRESETDONE),  
    .RESETEXCEPTION                     (),

    //----------------------------------------------------------------------------------------------
    //  PCIe Ports
    //----------------------------------------------------------------------------------------------
    .PCIERSTIDLE                        (GT_PCIERSTIDLE),        
    .PCIERSTTXSYNCSTART                 (GT_PCIERSTTXSYNCSTART), 
    .PCIEEQRXEQADAPTDONE                (GT_PCIEEQRXEQADAPTDONE),
    .PCIEUSERRATEDONE                   (GT_PCIEUSERRATEDONE),
             
    .PCIEUSERPHYSTATUSRST               (GT_PCIEUSERPHYSTATUSRST),    
    .PCIERATEQPLLPD                     (GT_PCIERATEQPLLPD),                    
    .PCIERATEQPLLRESET                  (GT_PCIERATEQPLLRESET),                 
    .PCIERATEIDLE                       (GT_PCIERATEIDLE),            
    .PCIESYNCTXSYNCDONE                 (GT_PCIESYNCTXSYNCDONE),                          
    .PCIERATEGEN3                       (pcierategen3),    
    .PCIEUSERGEN3RDY                    (GT_PCIEUSERGEN3RDY),   
    .PCIEUSERRATESTART                  (GT_PCIEUSERRATESTART),    
           
    //----------------------------------------------------------------------------------------------
    //  Serial Line Ports
    //----------------------------------------------------------------------------------------------
    .GTHRXP                             (GT_RXP),                                                   
    .GTHRXN                             (GT_RXN),   
   
    .GTHTXP                             (GT_TXP),                                                 
    .GTHTXN                             (GT_TXN),   

    //----------------------------------------------------------------------------------------------
    //  TX Data Ports
    //----------------------------------------------------------------------------------------------
    .TXDATA                             (txdata),                                     
    .TXCTRL0                            (txctrl0),
    .TXCTRL1                            (txctrl1),  
    .TXCTRL2                            (txctrl2),
    .TXDATAEXTENDRSVD                   ( 8'd0),                                

    //----------------------------------------------------------------------------------------------
    //  RX Data Ports
    //----------------------------------------------------------------------------------------------
    .RXDATA                             (rxdata),                                                    
    .RXCTRL0                            (rxctrl0),   
    .RXCTRL1                            (), 
    .RXCTRL2                            (),
    .RXCTRL3                            (), 
    .RXDATAEXTENDRSVD                   (),                                     
 
    //----------------------------------------------------------------------------------------------
    //  PHY Command Ports
    //----------------------------------------------------------------------------------------------
    .TXDETECTRX                         (GT_TXDETECTRX),                                            
    .TXELECIDLE                         (GT_TXELECIDLE),                                      
    .TXPDELECIDLEMODE                   ( 1'd0),                                                                                 
    .RXELECIDLEMODE                     ( 2'd0),                                
    .SIGVALIDCLK                        ( 1'd0),                                                                                    
    .TXPOLARITY                         ( 1'd0),                                              
    .RXPOLARITY                         (GT_RXPOLARITY),                                
    .TXPD                               (GT_POWERDOWN),                                           
    .RXPD                               (GT_POWERDOWN),                                           
    .TXRATE                             ({1'd0, GT_RATE}),                                                
    .RXRATE                             ({1'd0, GT_RATE}),                                                
    .TXRATEMODE                         ( 1'd0),                                                    
    .RXRATEMODE                         ( 1'd0),                                                    
 
    //----------------------------------------------------------------------------------------------
    //  PHY Status Ports
    //----------------------------------------------------------------------------------------------
    .RXVALID                            (GT_RXVALID),                                              
    .PHYSTATUS                          (GT_PHYSTATUS),                                            
    .RXELECIDLE                         (rxelecidle_int),                                           
    .RXSTATUS                           (GT_RXSTATUS),                                             
    .TXRATEDONE                         (),                                           
    .RXRATEDONE                         (GT_RXRATEDONE),                  
 
    //----------------------------------------------------------------------------------------------
    //  TX Driver Ports
    //----------------------------------------------------------------------------------------------
    .TXMARGIN                           (GT_TXMARGIN),                                           
    .TXSWING                            (GT_TXSWING),                                            
    .TXDEEMPH                           (GT_TXDEEMPH),                                                                     
    .TXDIFFCTRL                         (5'h14), //( 5'b11111), 
    .TXINHIBIT                          ( 1'd0),                                                  

    //----------------------------------------------------------------------------------------------
    //  TX Driver Ports (Gen3)
    //----------------------------------------------------------------------------------------------
    .TXPRECURSOR                        (GT_TXPRECURSOR),                                          
    .TXMAINCURSOR                       (GT_TXMAINCURSOR),                                         
    .TXPOSTCURSOR                       (GT_TXPOSTCURSOR),                                                                                     

    //----------------------------------------------------------------------------------------------
    //  PCS Reserved Ports
    //---------------------------------------------------------------------------------------------- 
    .PCSRSVDIN                          (16'h0001),                             // CHECK                                                                               
    .PCSRSVDOUT                         (pcsrsvdout),     
    
    //----------------------------------------------------------------------------------------------
    //  RX Monitor Ports
    //----------------------------------------------------------------------------------------------
    .RXMONITORSEL                       ( 2'd0), 
    .RXMONITOROUT                       (),                                                                                                                                                                                                            
                                                                 
    //----------------------------------------------------------------------------------------------
    //  Comma Detect & Align Ports
    //----------------------------------------------------------------------------------------------
    .RXCOMMADETEN                       ( 1'd1),                  
    .RXMCOMMAALIGNEN                    (!pcierategen3),          
    .RXPCOMMAALIGNEN                    (!pcierategen3),          
                                                                                 
    .RXCOMMADET                         (),                                            
    .RXBYTEISALIGNED                    (),                                        
    .RXBYTEREALIGN                      (),                                                                                                                 
                                                                                                    
    //----------------------------------------------------------------------------------------------
    // 8B10B Ports
    //----------------------------------------------------------------------------------------------
    .TX8B10BBYPASS                      ( 8'd0),                                                  
    .TX8B10BEN                          (!pcierategen3),                            
    .RX8B10BEN                          (!pcierategen3),                            
           
    //----------------------------------------------------------------------------------------------
    //  TX Buffer Ports
    //----------------------------------------------------------------------------------------------
    .TXBUFSTATUS                        (),                                                        
                                                                                                    
    //----------------------------------------------------------------------------------------------
    //  RX Buffer Ports
    //----------------------------------------------------------------------------------------------
    .RXBUFRESET                         (GT_RXBUFRESET),                                          
    .RXBUFSTATUS                        (),                
                      
    //----------------------------------------------------------------------------------------------
    //  Clock Correction Ports
    //----------------------------------------------------------------------------------------------
    .RXCLKCORCNT                        (),                            
                    
    //----------------------------------------------------------------------------------------------
    //  Channel Bonding Ports (disable)
    //----------------------------------------------------------------------------------------------
    .RXCHBONDEN                         ( 1'd0),                                         
    .RXCHBONDI                          ( 5'd0),                                         
    .RXCHBONDLEVEL                      ( 3'd0),                                         
    .RXCHBONDMASTER                     ( 1'd0),                                         
    .RXCHBONDSLAVE                      ( 1'd0),                                         
                                                                                    
    .RXCHANBONDSEQ                      (),                                         
    .RXCHANISALIGNED                    (),                                         
    .RXCHANREALIGN                      (),                                         
    .RXCHBONDO                          (),                                                                                                                                                                       
 
    //----------------------------------------------------------------------------------------------
    //  TX Phase Alignment Ports
    //----------------------------------------------------------------------------------------------
    .TXPHALIGN                          ( 1'd0),
    .TXPHALIGNEN                        ( 1'd0),
    .TXPHDLYPD                          ( 1'd0),
    .TXPHDLYRESET                       ( 1'd0),
    .TXPHDLYTSTCLK                      ( 1'd0),
    .TXPHINIT                           ( 1'd0),
    .TXPHOVRDEN                         ( 1'd0),
   
    .TXPHALIGNDONE                      (GT_TXPHALIGNDONE),
    .TXPHINITDONE                       (),
   
    //----------------------------------------------------------------------------------------------
    //  TX Delay Alignment Ports
    //----------------------------------------------------------------------------------------------
    .TXDLYBYPASS                        ( 1'd0),
    .TXDLYEN                            ( 1'd0),
    .TXDLYHOLD                          ( 1'd0),
    .TXDLYOVRDEN                        ( 1'd0),
    .TXDLYSRESET                        ( 1'd0),
    .TXDLYUPDOWN                        ( 1'd0),
       
    .TXDLYSRESETDONE                    (),       
          
    //----------------------------------------------------------------------------------------------
    //  TX Auto Sync Alignment Ports 
    //----------------------------------------------------------------------------------------------
    .TXSYNCALLIN                        (GT_TXSYNCALLIN),
    .TXSYNCIN                           (GT_TXSYNCIN),
    .TXSYNCMODE                         (MASTER_LANE),                                         
                
    .TXSYNCDONE                         (),
    .TXSYNCOUT                          (GT_TXSYNCOUT),

    //----------------------------------------------------------------------------------------------
    //  RX Phase Alignment Ports (disable)
    //----------------------------------------------------------------------------------------------
    .RXPHALIGN                          ( 1'd0),
    .RXPHALIGNEN                        ( 1'd0),
    .RXPHDLYPD                          ( 1'd0),
    .RXPHDLYRESET                       ( 1'd0),
    .RXPHOVRDEN                         ( 1'd0),
   
    .RXPHALIGNDONE                      (),
    .RXPHALIGNERR                       (),
       
    //----------------------------------------------------------------------------------------------
    //  RX Delay Alignment Ports (disable)
    //----------------------------------------------------------------------------------------------
    .RXDLYBYPASS                        ( 1'd1),
    .RXDLYEN                            ( 1'd0),
    .RXDLYOVRDEN                        ( 1'd0),
    .RXDLYSRESET                        ( 1'd0),
   
    .RXDLYSRESETDONE                    (),                                           
        
    //----------------------------------------------------------------------------------------------
    //  RX Auto Sync Alignment Ports (disable)
    //----------------------------------------------------------------------------------------------
    .RXSYNCALLIN                        ( 1'd0),
    .RXSYNCIN                           ( 1'd0),
    .RXSYNCMODE                         ( 1'd0),                                                    
                                                                                                    
    .RXSYNCDONE                         (),                                                
    .RXSYNCOUT                          (),    
       
    //----------------------------------------------------------------------------------------------
    //  Gearbox Ports 
    //----------------------------------------------------------------------------------------------
    .TXHEADER                           ( 6'd0), 
    .TXLATCLK                           ( 1'd0),                                                    
    .TXSEQUENCE                         ( 7'd0),                                                    
    .RXGEARBOXSLIP                      ( 1'd0),  
    .RXLATCLK                           ( 1'd0),  
    .RXSLIDE                            ( 1'd0),                                                    
                                                                                                    
    .RXDATAVALID                        (),                 
    .RXHEADER                           (),                                                         
    .RXHEADERVALID                      (), 
    .RXSLIDERDY                         (),                                                         
    .RXSTARTOFSEQ                       (),                             
                   
    //----------------------------------------------------------------------------------------------
    //  RX Slip Ports 
    //----------------------------------------------------------------------------------------------
    .RXSLIPOUTCLK                       ( 1'd0),
    .RXSLIPPMA                          ( 1'd0),   
                                                                   
    .RXSLIPDONE                         (),     
    .RXSLIPOUTCLKRDY                    (),
    .RXSLIPPMARDY                       (),             
       
    //----------------------------------------------------------------------------------------------
    //  RX LPM Ports 
    //----------------------------------------------------------------------------------------------
    .RXLPMEN                            (!pcierategen3),    
    .RXLPMGCHOLD                        ( 1'b0),            
    .RXLPMGCOVRDEN                      ( 1'b0),
    .RXLPMHFHOLD                        ( 1'b0),            
    .RXLPMHFOVRDEN                      ( 1'b0),
    .RXLPMLFHOLD                        ( 1'b0),         
    .RXLPMLFKLOVRDEN                    ( 1'b0), 
    .RXLPMOSHOLD                        ( 1'b0),            
    .RXLPMOSOVRDEN                      ( 1'b0),
                                                                                                    
    //----------------------------------------------------------------------------------------------
    //  RX DFE Ports
    //----------------------------------------------------------------------------------------------
    .RXDFEAGCCTRL                       ( 2'h1), //( 2'b00),   
    .RXDFEAGCHOLD                       ( 1'b0),            
    .RXDFEAGCOVRDEN                     ( 1'b0),
    .RXDFECFOKFCNUM                     ( 4'b0000),                             
    .RXDFECFOKFEN                       ( 1'b0),                                
    .RXDFECFOKFPULSE                    ( 1'b0),                                
    .RXDFECFOKHOLD                      ( 1'b0),                                
    .RXDFECFOKOVREN                     ( 1'b0),                                
    .RXDFEKHHOLD                        ( 1'b0),
    .RXDFEKHOVRDEN                      ( 1'b0),
    .RXDFELFHOLD                        ( 1'b0),          
    .RXDFELFOVRDEN                      ( 1'b0),
    .RXDFELPMRESET                      (GT_RXDFELPMRESET),
    .RXDFETAP2HOLD                      ( 1'b0),
    .RXDFETAP2OVRDEN                    ( 1'b0),
    .RXDFETAP3HOLD                      ( 1'b0),
    .RXDFETAP3OVRDEN                    ( 1'b0),
    .RXDFETAP4HOLD                      ( 1'b0),
    .RXDFETAP4OVRDEN                    ( 1'b0),
    .RXDFETAP5HOLD                      ( 1'b0),
    .RXDFETAP5OVRDEN                    ( 1'b0),
    .RXDFETAP6HOLD                      ( 1'b0),
    .RXDFETAP6OVRDEN                    ( 1'b0),
    .RXDFETAP7HOLD                      ( 1'b0),
    .RXDFETAP7OVRDEN                    ( 1'b0),
    .RXDFETAP8HOLD                      ( 1'b0),
    .RXDFETAP8OVRDEN                    ( 1'b0),
    .RXDFETAP9HOLD                      ( 1'b0),
    .RXDFETAP9OVRDEN                    ( 1'b0),
    .RXDFETAP10HOLD                     ( 1'b0),
    .RXDFETAP10OVRDEN                   ( 1'b0),
    .RXDFETAP11HOLD                     ( 1'b0),
    .RXDFETAP11OVRDEN                   ( 1'b0),
    .RXDFETAP12HOLD                     ( 1'b0),
    .RXDFETAP12OVRDEN                   ( 1'b0),
    .RXDFETAP13HOLD                     ( 1'b0),
    .RXDFETAP13OVRDEN                   ( 1'b0),
    .RXDFETAP14HOLD                     ( 1'b0),
    .RXDFETAP14OVRDEN                   ( 1'b0),
    .RXDFETAP15HOLD                     ( 1'b0),
    .RXDFETAP15OVRDEN                   ( 1'b0),
    .RXDFEUTHOLD                        ( 1'b0),
    .RXDFEUTOVRDEN                      ( 1'b0),
    .RXDFEVPHOLD                        ( 1'b0),
    .RXDFEVPOVRDEN                      ( 1'b0),
    .RXDFEXYDEN                         ( 1'b1),                                                                                                    
    
    //----------------------------------------------------------------------------------------------
    //  TX PI Ports
    //----------------------------------------------------------------------------------------------
    .TXPIPPMEN                          ( 1'd0),
    .TXPIPPMOVRDEN                      ( 1'd0),
    .TXPIPPMPD                          ( 1'd0),
    .TXPIPPMSEL                         ( 1'd0),
    .TXPIPPMSTEPSIZE                    ( 5'd0),
    .TXPISOPD                           ( 1'd0),   
    
    //----------------------------------------------------------------------------------------------
    //  RX CDR Ports
    //----------------------------------------------------------------------------------------------
    .CDRSTEPDIR                         ( 1'b0),                                 
    .CDRSTEPSQ                          ( 1'b0),                                
    .CDRSTEPSX                          ( 1'b0),                               
    .RXCDRFREQRESET                     (GT_RXCDRFREQRESET),   //*****
    .RXCDRHOLD                          (GT_RXCDRHOLD),
    .RXCDROVRDEN                        ( 1'd0),
    .RXCDRRESET                         (rxcdrreset_int),
    
    .RXCDRLOCK                          (GT_RXCDRLOCK),    
    .RXCDRPHDONE                        (), 
       
    //----------------------------------------------------------------------------------------------
    //  Eye Scan Ports
    //----------------------------------------------------------------------------------------------                                          
    .EYESCANRESET                       ( 1'd0),                                             
    .EYESCANTRIGGER                     ( 1'd0),                                             
                                                                                            
    .EYESCANDATAERROR                   (),           
       
    //----------------------------------------------------------------------------------------------
    //  RX OS Ports
    //----------------------------------------------------------------------------------------------
    .RXOSCALRESET                       ( 1'b0),
    .RXOSHOLD                           ( 1'b0),
    .RXOSOVRDEN                         ( 1'b0),    
 
    .RXOSINTDONE                        (),                                                         
    .RXOSINTSTARTED                     (),                                                         
    .RXOSINTSTROBEDONE                  (),                                                         
    .RXOSINTSTROBESTARTED               (),         
           
    //----------------------------------------------------------------------------------------------
    //  DRP Ports
    //----------------------------------------------------------------------------------------------
    .DRPCLK                             (GT_DRPCLK), 
    .DRPRST                             ( 1'd0),                                                                                
    .DRPADDR                            (GT_DRPADDR),                                                    
    .DRPEN                              (GT_DRPEN),                                                    
    .DRPWE                              (GT_DRPWE), 
    .DRPDI                              (GT_DRPDI),                                                    
        
    .DRPRDY                             (GT_DRPRDY),                                                         
    .DRPDO                              (GT_DRPDO),                      
 
    //----------------------------------------------------------------------------------------------
    //  Loopback & PRBS Ports
    //----------------------------------------------------------------------------------------------
    .LOOPBACK                           (GT_LOOPBACK),      
    .TXPRBSSEL                          (GT_PRBSSEL),                                                    
    .RXPRBSSEL                          (GT_PRBSSEL),  
    .TXPRBSFORCEERR                     (GT_TXPRBSFORCEERR),  
    .RXPRBSCNTRESET                     (GT_RXPRBSCNTRESET),  
                   
    .RXPRBSERR                          (GT_RXPRBSERR),                                                
    .RXPRBSLOCKED                       (GT_RXPRBSLOCKED),       

    //----------------------------------------------------------------------------------------------
    //  Digital Monitor Ports                                                                             
    //----------------------------------------------------------------------------------------------
    .DMONFIFORESET                      ( 1'd0),                                                    
    .DMONITORCLK                        ( 1'd0),                                                    
    
    .DMONITOROUT                        (),    
    .DMONITOROUTCLK                     (),                                             
      
    //----------------------------------------------------------------------------------------------
    //  USB Ports
    //----------------------------------------------------------------------------------------------
    .TXONESZEROS                        (GT_TXONESZEROS),
    .RXEQTRAINING                       (GT_RXEQTRAINING),
    .RXTERMINATION                      (GT_RXTERMINATION),    
    
    .POWERPRESENT                       (GT_POWERPRESENT),           
        
    //----------------------------------------------------------------------------------------------
    //  USB LFPS Ports
    //----------------------------------------------------------------------------------------------
    .TXLFPSTRESET                       ( 1'b0),      
    .TXLFPSU2LPEXIT                     ( 1'b0),
    .TXLFPSU3WAKE                       ( 1'b0),
    
    .RXLFPSTRESETDET                    (),             
    .RXLFPSU2LPEXITDET                  (),             
    .RXLFPSU3WAKEDET                    (),            
      
    //----------------------------------------------------------------------------------------------
    //  SATA Ports 
    //----------------------------------------------------------------------------------------------
    .TXCOMINIT                          ( 1'd0),                                                    
    .TXCOMSAS                           ( 1'd0),                                                    
    .TXCOMWAKE                          ( 1'd0),                                                    

    .TXCOMFINISH                        (),                                                         
    .RXCOMINITDET                       (),                                                         
    .RXCOMSASDET                        (),                                                         
    .RXCOMWAKEDET                       (),                                                    

    //----------------------------------------------------------------------------------------------
    //  QPI
    //----------------------------------------------------------------------------------------------
    .RXQPIEN                            ( 1'd0),
    .TXQPIBIASEN                        ( 1'b0),                                
    .TXQPIWEAKPUP                       ( 1'b0),                              
    
    .RXQPISENN                          (),
    .RXQPISENP                          (),
    .TXQPISENN                          (),
    .TXQPISENP                          (),

    //----------------------------------------------------------------------------------------------
    //  GT Ports
    //----------------------------------------------------------------------------------------------
    .FREQOS                             ( 1'd0),    
    .GTRSVD                             (16'd0),
    .INCPCTRL                           ( 1'd0),
    .RXAFECFOKEN                        ( 1'd0),                                
    .RXCKCALRESET                       ( 1'b0),                                
    .RXCKCALSTART                       ( 7'd0),                                
    .TSTIN                              (20'h00000),                                                
    .TXDCCFORCESTART                    ( 1'b0),                                
    .TXDCCRESET                         ( 1'b0),                                
    .TXMUXDCDEXHOLD                     ( 1'b0),                                
    .TXMUXDCDORWREN                     ( 1'b0),                                
                                                                                   
    .PINRSRVDAS                         (),                                     
    .RXCKCALDONE                        (),                                     
    .TXDCCDONE                          ()                                      
);

end
endgenerate


//--------------------------------------------------------------------------------------------------
//  Input Port Remapping
//--------------------------------------------------------------------------------------------------    
assign txdata[ 63: 0] = GT_TXDATA;
assign txdata[127:64] = 64'd0;

assign txctrl0[ 1:0] = 2'd0;
assign txctrl0[   2] = GT_TXDATA_VALID;
assign txctrl0[   3] = GT_TXSTART_BLOCK;
assign txctrl0[ 5:4] = GT_TXSYNC_HEADER;
assign txctrl0[15:6] = 10'd0;

assign txctrl1[   0] = GT_TXCOMPLIANCE;
assign txctrl1[15:1] = 15'd0;

assign txctrl2[ 1:0] = GT_TXDATAK;
assign txctrl2[ 7:2] = 6'd0;



//--------------------------------------------------------------------------------------------------
//  GT Channel Outputs
//--------------------------------------------------------------------------------------------------
assign GT_RXDATA         = rxdata[63:0];

assign GT_RXDATAK        = rxctrl0[1:0];
assign GT_RXDATA_VALID   = rxctrl0[2];
assign GT_RXSTART_BLOCK  = {rxctrl0[6], rxctrl0[3]};
assign GT_RXSYNC_HEADER  = rxctrl0[5:4];
assign GT_GEN34_EIOS_DET = rxctrl0[7]; 

assign GT_PCIERATEGEN3   = pcierategen3;
assign GT_QPLLRATE       = pcsrsvdout[2:0];

assign GT_RXELECIDLE = rxelecidle_int;


endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_gt_gt_common.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
//  Design :  PHY Wrapper
//  Module :  GT Common
//--------------------------------------------------------------------------------------------------

`timescale 1ps / 1ps

//--------------------------------------------------------------------------------------------------
//  GT Common Module
//--------------------------------------------------------------------------------------------------
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_gt_gt_common #
(
    parameter         PHY_SIM_EN      = "FALSE",
    parameter         PHY_GT_XCVR     = "GTY",
    parameter integer PHY_MAX_SPEED   = 4,
    parameter integer PHY_REFCLK_FREQ = 0    
)
(    
    //----------------------------------------------------------------------------------------------
    //  Clock Ports
    //----------------------------------------------------------------------------------------------
    input                               GTCOM_REFCLK,
    
    output                              GTCOM_QPLL0OUTCLK,
    output                              GTCOM_QPLL0OUTREFCLK,
    output                              GTCOM_QPLL0LOCK,
    
    output                              GTCOM_QPLL1OUTCLK,
    output                              GTCOM_QPLL1OUTREFCLK,
    output                              GTCOM_QPLL1LOCK,
    
    //----------------------------------------------------------------------------------------------
    //  Reset Ports
    //----------------------------------------------------------------------------------------------
    input                               GTCOM_QPLL0PD,
    input                               GTCOM_QPLL0RESET, 
 
    input                               GTCOM_QPLL1PD,
    input                               GTCOM_QPLL1RESET,
            
    //----------------------------------------------------------------------------------------------
    //  PCIe Ports
    //----------------------------------------------------------------------------------------------
    input       [ 2:0]                  GTCOM_QPLLRATE,
    
    //----------------------------------------------------------------------------------------------
    //  DRP Ports
    //----------------------------------------------------------------------------------------------
    input                               GTCOM_DRPCLK,                                        
    input       [15:0]                  GTCOM_DRPADDR,                                       
    input                               GTCOM_DRPEN,                                             
    input                               GTCOM_DRPWE,     
    input       [15:0]                  GTCOM_DRPDI,                                      
                                                                
    output                              GTCOM_DRPRDY,    
    output      [15:0]                  GTCOM_DRPDO
);                                                      
    
    //----------------------------------------------------------------------------------------------
    //  QPLL[0/1]_FBDIV - QPLL Feedback (N) Divider (Gen1/Gen2)
    //----------------------------------------------------------------------------------------------
    localparam [ 7:0] QPLL_FBDIV = (PHY_REFCLK_FREQ == 2) ? 8'd40 : 
                                   (PHY_REFCLK_FREQ == 1) ? 8'd80 : 8'd100;
    
    
    
    //----------------------------------------------------------------------------------------------
    //  QPLL[1/0]_FBDIV_G34 - QPLL Feedback (N) Divider (Gen3/Gen4)
    //----------------------------------------------------------------------------------------------    
    localparam [ 7:0] QPLL_FBDIV_G3 = (PHY_REFCLK_FREQ == 2) ? 8'd32  : 
                                      (PHY_REFCLK_FREQ == 1) ? 8'd64  : 8'd80;
    
    localparam [ 7:0] QPLL_FBDIV_G4 = (PHY_REFCLK_FREQ == 2) ? 8'd64  : 
                                      (PHY_REFCLK_FREQ == 1) ? 8'd128 : 8'd160;
    
    localparam [ 7:0] QPLL_FBDIV_G34 = (PHY_MAX_SPEED == 4) ? QPLL_FBDIV_G4 : QPLL_FBDIV_G3;



    //----------------------------------------------------------------------------------------------
    //  QPLL[1/0]_CFG2_G3 - QPLL Configuration (Gen3 and Gen4)
    //    [6] : 1'b0 = Select upper band VCO
    //        : 1'b1 = Select lower band VCO
    //----------------------------------------------------------------------------------------------  
    localparam [15:0] QPLL_CFG2_G3 = (PHY_MAX_SPEED == 4) ? 16'h0000 : 16'h0040;



//--------------------------------------------------------------------------------------------------
//  GTY Common
//--------------------------------------------------------------------------------------------------    

generate
  if (PHY_GT_XCVR == "GTY" || PHY_GT_XCVR == "GTY64") begin: GTY_CHANNEL
//--------------------------------------------------------------------------------------------------
//  GTY Common
//--------------------------------------------------------------------------------------------------
GTYE4_COMMON #
(   
    //---------------------------------------------------------------------------------------------- 
    //  Simulation Attributes
    //----------------------------------------------------------------------------------------------      
    .SIM_MODE                           ("FAST"),                                                                                                                                                                                      
    .SIM_RESET_SPEEDUP                  ("TRUE"),                                                                                              
    //.SIM_VERSION                        (1),                                                                          

    //----------------------------------------------------------------------------------------------               
    //  Clock Attributes
    //----------------------------------------------------------------------------------------------    
    .RXRECCLKOUT0_SEL                   ( 2'b00),
    .RXRECCLKOUT1_SEL                   ( 2'b00),                    

    //----------------------------------------------------------------------------------------------
    //  QPLL0 Attributes 
    //----------------------------------------------------------------------------------------------    
    .AEN_QPLL0_FBDIV                    (1'b1),                                 
    .QPLL0CLKOUT_RATE                   ("HALF"),                              
    .QPLL0_CFG0                         (16'h001D),                             
    .QPLL0_CFG1                         (16'h0000),                             
    .QPLL0_CFG1_G3                      (16'h0000),                             
    .QPLL0_CFG2                         (16'h0040),                             
    .QPLL0_CFG2_G3                      (QPLL_CFG2_G3),                        
    .QPLL0_CFG3                         (16'h0120),                  
    .QPLL0_CFG4                         (16'h0000),
    .QPLL0_CP                           (10'b0000011111),                       // Optimized for PCIe PLL compliance
    .QPLL0_CP_G3                        (10'b0000011111),                       // Optimized for PCIe PLL compliance
    .QPLL0_FBDIV                        (QPLL_FBDIV),
    .QPLL0_FBDIV_G3                     (QPLL_FBDIV_G34),
    .QPLL0_INIT_CFG0                    (16'b0000000000000000),
    .QPLL0_INIT_CFG1                    ( 8'b00000000),
    .QPLL0_LOCK_CFG                     (16'h05FC),                             // [10] : 1'b1 = Auto VCO
    .QPLL0_LOCK_CFG_G3                  (16'h05FC),                             // [10] : 1'b1 = Auto VCO
    .QPLL0_LPF                          (10'b0000010101),                       // Optimized for PCIe PLL compliance
    .QPLL0_LPF_G3                       (10'b0000010101),                       // Optimized for PCIe PLL compliance
    .QPLL0_PCI_EN                       ( 1'b1),                                
    .QPLL0_RATE_SW_USE_DRP              ( 1'b0),                                // Advance PCIe feature
    .QPLL0_REFCLK_DIV                   (1),
    .QPLL0_SDM_CFG0                     (16'b0000000011000000),                
    .QPLL0_SDM_CFG1                     (16'b0000000000000000),
    .QPLL0_SDM_CFG2                     (16'b0000000000000000),
                     
    //---------------------------------------------------------------------------------------------- 
    //  QPLL1 Attributes               
    //----------------------------------------------------------------------------------------------    
    .AEN_QPLL1_FBDIV                    (1'b1),                                 
    .QPLL1CLKOUT_RATE                   ("HALF"),                              
    .QPLL1_CFG0                         (16'h001D),                             
    .QPLL1_CFG1                         (16'h0000),                             
    .QPLL1_CFG1_G3                      (16'h0000),                             
    .QPLL1_CFG2                         (16'h0040),                             
    .QPLL1_CFG2_G3                      (QPLL_CFG2_G3),                         
    .QPLL1_CFG3                         (16'h0120),                  
    .QPLL1_CFG4                         (16'h0000),
    .QPLL1_CP                           (10'b0000011111),                       // Optimized for PCIe PLL compliance
    .QPLL1_CP_G3                        (10'b0000011111),                       // Optimized for PCIe PLL compliance
    .QPLL1_FBDIV                        (QPLL_FBDIV),
    .QPLL1_FBDIV_G3                     (QPLL_FBDIV_G34),
    .QPLL1_INIT_CFG0                    (16'b0000000000000000),
    .QPLL1_INIT_CFG1                    ( 8'b00000000),
    .QPLL1_LOCK_CFG                     (16'h05FC),                             // [10] : 1'b1 = Auto VCO
    .QPLL1_LOCK_CFG_G3                  (16'h05FC),                             // [10] : 1'b1 = Auto VCO
    .QPLL1_LPF                          (10'b0000010101),                       // Optimized for PCIe PLL compliance
    .QPLL1_LPF_G3                       (10'b0000010101),                       // Optimized for PCIe PLL compliance
    .QPLL1_PCI_EN                       ( 1'b1),                               
    .QPLL1_RATE_SW_USE_DRP              ( 1'b0),                                // Advance PCIe feature
    .QPLL1_REFCLK_DIV                   (1),
    .QPLL1_SDM_CFG0                     (16'b0000000011000000),                 
    .QPLL1_SDM_CFG1                     (16'b0000000000000000),
    .QPLL1_SDM_CFG2                     (16'b0000000000000000),
 
    //----------------------------------------------------------------------------------------------
    //  PPF Attributes                                                         
    //----------------------------------------------------------------------------------------------      
    .PPF0_CFG                           (16'h0FFF),                            
    .PPF1_CFG                           (16'h0FFF),                           
    
    //----------------------------------------------------------------------------------------------
    //  Bias Attributes                                                          
    //----------------------------------------------------------------------------------------------
    .BIAS_CFG0                          (16'b0000000000000000),
    .BIAS_CFG1                          (16'b0000000000000000),
    .BIAS_CFG2                          (16'b0011000000000000),                 // Optimized for PCIe PLL compliance
    .BIAS_CFG3                          (16'b0000000001000000),                 
    .BIAS_CFG4                          (16'b0000000000000000),    
    .BIAS_CFG_RSVD                      (10'b0000000000),  
       
    //---------------------------------------------------------------------------------------------- 
    //  SDM0 Attributes                                                          
    //----------------------------------------------------------------------------------------------
    .A_SDM0TOGGLE                       ( 1'b0),
    .AEN_SDM0TOGGLE                     ( 1'b0),
    .SDM0INITSEED0_0                    (16'b0000000000000000),
    .SDM0INITSEED0_1                    ( 9'b000000000),
    
    //---------------------------------------------------------------------------------------------- 
    //  SDM1 Attributes                                                          
    //----------------------------------------------------------------------------------------------     
    .A_SDM1DATA_HIGH                    ( 9'b000000000),
    .A_SDM1DATA_LOW                     (16'b0000000000000000),
    .A_SDM1TOGGLE                       ( 1'b0),
    .AEN_SDM1TOGGLE                     ( 1'b0),
    .SDM1INITSEED0_0                    (16'b0000000000000000),
    .SDM1INITSEED0_1                    ( 9'b000000000),     
          
    //----------------------------------------------------------------------------------------------
    //  Reserved & MISC Attributes                                                         
    //----------------------------------------------------------------------------------------------            
    .COMMON_CFG0                        (16'b0000000000000000),
    .COMMON_CFG1                        (16'b0000000000000000),
    .POR_CFG                            (16'b0000000000001011),                 // CHECK      
    .RSVD_ATTR0                         (16'b0000000000000001),                 // CHECK
    .RSVD_ATTR1                         (16'b0000000000000000),    
    .RSVD_ATTR2                         (16'b0000000000000001),                 // CHECK                
    .RSVD_ATTR3                         (16'b0000000000000000),
    .SARC_ENB                           ( 1'b0),
    .SARC_SEL                           ( 1'b0),

    //----------------------------------------------------------------------------------------------
    //  MicroBlaze Attributes                                                         
    //----------------------------------------------------------------------------------------------
    .UB_CFG0                            (16'h0),
    .UB_CFG1                            (16'h0),
    .UB_CFG2                            (16'h0),
    .UB_CFG3                            (16'h0),
    .UB_CFG4                            (16'h0),
    .UB_CFG5                            (16'h0),
    .UB_CFG6                            (16'h0)
)
gtye4_common_smsw_i 
(       
    //----------------------------------------------------------------------------------------------
    //  QPLL0 Clock Ports
    //----------------------------------------------------------------------------------------------
    .GTGREFCLK0                         ( 1'd0), 
    .GTREFCLK00                         (GTCOM_REFCLK),                         
    .GTREFCLK10                         ( 1'd0),
    .GTNORTHREFCLK00                    ( 1'd0),
    .GTNORTHREFCLK10                    ( 1'd0),
    .GTSOUTHREFCLK00                    ( 1'd0),
    .GTSOUTHREFCLK10                    ( 1'd0),
   
    .REFCLKOUTMONITOR0                  (),
    .RXRECCLK0SEL                       (),
    
    //----------------------------------------------------------------------------------------------
    //  QPLL1 Clock Ports
    //----------------------------------------------------------------------------------------------
    .GTGREFCLK1                         ( 1'd0),
    .GTREFCLK01                         (GTCOM_REFCLK),
    .GTREFCLK11                         ( 1'd0),
    .GTNORTHREFCLK01                    ( 1'd0),    
    .GTNORTHREFCLK11                    ( 1'd0),
    .GTSOUTHREFCLK01                    ( 1'd0),
    .GTSOUTHREFCLK11                    ( 1'd0),        
        
    .REFCLKOUTMONITOR1                  (),  
    .RXRECCLK1SEL	                      (), 
        
    //----------------------------------------------------------------------------------------------
    //  QPLL0 Ports
    //----------------------------------------------------------------------------------------------
    .QPLL0CLKRSVD0                      ( 1'd0),
    .QPLL0CLKRSVD1                      ( 1'd0),                              
    .QPLL0FBDIV                         ( 8'd0),                                // CHECK
    .QPLL0LOCKDETCLK                    ( 1'd0),
    .QPLL0LOCKEN                        ( 1'd1),
    .QPLL0PD                            (GTCOM_QPLL0PD),                        
    .QPLL0REFCLKSEL                     ( 3'd1),                                                          
    .QPLL0RESET                         (GTCOM_QPLL0RESET),                     
       
    .QPLL0FBCLKLOST                     (),
    .QPLL0LOCK                          (GTCOM_QPLL0LOCK),
    .QPLL0OUTCLK                        (GTCOM_QPLL0OUTCLK),
    .QPLL0OUTREFCLK                     (GTCOM_QPLL0OUTREFCLK),
    .QPLL0REFCLKLOST                    (),     
    .QPLLDMONITOR0                      (),                                                                      
                                               
    //----------------------------------------------------------------------------------------------
    //  QPLL1 Ports
    //----------------------------------------------------------------------------------------------
    .QPLL1CLKRSVD0                      ( 1'd0),
    .QPLL1CLKRSVD1                      ( 1'd0),                                
    .QPLL1FBDIV                         ( 8'd0),                                // CHECK
    .QPLL1LOCKDETCLK                    ( 1'd0),
    .QPLL1LOCKEN                        ( 1'd1),
    .QPLL1PD                            (GTCOM_QPLL1PD),
    .QPLL1REFCLKSEL                     ( 3'd1),                        
    .QPLL1RESET                         (GTCOM_QPLL1RESET),      
     
    .QPLL1FBCLKLOST                     (),  
    .QPLL1LOCK                          (GTCOM_QPLL1LOCK),       
    .QPLL1OUTCLK                        (GTCOM_QPLL1OUTCLK),     
    .QPLL1OUTREFCLK                     (GTCOM_QPLL1OUTREFCLK),                       
    .QPLL1REFCLKLOST                    (),  
    .QPLLDMONITOR1                      (),            
         
    //----------------------------------------------------------------------------------------------
    //  PCIe Ports
    //----------------------------------------------------------------------------------------------
    .PCIERATEQPLL0                      (GTCOM_QPLLRATE),           
    .PCIERATEQPLL1                      (GTCOM_QPLLRATE),       
                                                                                                       
    //----------------------------------------------------------------------------------------------
    //  DRP Ports
    //----------------------------------------------------------------------------------------------
    .DRPCLK                             (GTCOM_DRPCLK),                                        
    .DRPADDR                            (GTCOM_DRPADDR),                                       
    .DRPEN                              (GTCOM_DRPEN),                                             
    .DRPWE                              (GTCOM_DRPWE),     
    .DRPDI                              (GTCOM_DRPDI),                                      
                                                                         
    .DRPRDY                             (GTCOM_DRPRDY),    
    .DRPDO                              (GTCOM_DRPDO),                                      
        
    //----------------------------------------------------------------------------------------------
    //  rCal Ports
    //----------------------------------------------------------------------------------------------        
    .RCALENB                            ( 1'd1),          
                                                                                                        
    //----------------------------------------------------------------------------------------------
    //  Band Gap Ports
    //----------------------------------------------------------------------------------------------
    .BGBYPASSB                          ( 1'b1),                                
    .BGMONITORENB                       ( 1'b1),                                
    .BGPDB                              ( 1'b1),  
    .BGRCALOVRD                         ( 5'b11111),                                 
    .BGRCALOVRDENB                      ( 1'b1),                                                            
        
    //----------------------------------------------------------------------------------------------
    //  SDM0 Ports
    //----------------------------------------------------------------------------------------------
    .SDM0DATA                           (25'd0),
    .SDM0RESET                          ( 1'd0),
    .SDM0TOGGLE                         ( 1'd0), 
    .SDM0WIDTH                          ( 2'd0),
    
    .SDM0FINALOUT                       (),
    .SDM0TESTDATA                       (),

    //----------------------------------------------------------------------------------------------
    //  SDM1 Ports
    //----------------------------------------------------------------------------------------------
    .SDM1DATA                           (25'd0),
    .SDM1RESET                          ( 1'd0),
    .SDM1TOGGLE                         ( 1'd0), 
    .SDM1WIDTH                          ( 2'd0),
    
    .SDM1FINALOUT                       (),
    .SDM1TESTDATA                       (),

    //----------------------------------------------------------------------------------------------
    //  TCON Ports
    //----------------------------------------------------------------------------------------------
    //.TCONGPI                            (10'd0),
    //.TCONPOWERUP                        ( 1'd0),
    //.TCONRESET                          ( 2'd0),
    //.TCONRSVDIN1                        ( 2'd0),
    
    //.TCONGPO                            (),
    //.TCONRSVDOUT0                       (),

    //----------------------------------------------------------------------------------------------
    //  Reserved & MISC Ports
    //----------------------------------------------------------------------------------------------
    .PMARSVD0                           ( 8'd0),            
    .PMARSVD1                           ( 8'd0),  
    .QPLLRSVD1                          ( 8'd0),
    .QPLLRSVD2                          ( 5'd0),               
    .QPLLRSVD3                          ( 5'd0),          
    .QPLLRSVD4                          ( 8'd0),                   

    .PMARSVDOUT0                        (),
    .PMARSVDOUT1                        (),

    //----------------------------------------------------------------------------------------------
    //  MicroBlaze Ports
    //----------------------------------------------------------------------------------------------
    .UBCFGSTREAMEN                      ( 1'b0),
    .UBDO                               ( 16'h0),
    .UBDRDY                             ( 1'b0),
    .UBENABLE                           ( 1'b0),
    .UBGPI                              ( 2'b0),
    .UBINTR                             ( 2'b0),
    .UBIOLMBRST                         ( 1'b0),
    .UBMBRST                            ( 1'b0),
    .UBMDMCAPTURE                       ( 1'b0),
    .UBMDMDBGRST                        ( 1'b0),
    .UBMDMDBGUPDATE                     ( 1'b0),
    .UBMDMREGEN                         ( 4'b0),
    .UBMDMSHIFT                         ( 1'b0),
    .UBMDMSYSRST                        ( 1'b0),
    .UBMDMTCK                           ( 1'b0),
    .UBMDMTDI                           ( 1'b0),

    .UBDADDR                            (),
    .UBDEN                              (),
    .UBDI                               (),
    .UBDWE                              (),
    .UBMDMTDO                           (),
    .UBRSVDOUT                          (),
    .UBTXUART                           ()

);

end else begin: GTH_COMMON
GTHE4_COMMON #
(   
    //---------------------------------------------------------------------------------------------- 
    //  Simulation Attributes
    //----------------------------------------------------------------------------------------------      
    .SIM_MODE                           ("FAST"),                                                                                                                                                                                      
    .SIM_RESET_SPEEDUP                  ("TRUE"),                                                                                              
    //.SIM_VERSION                        (1),                                                                          

    //----------------------------------------------------------------------------------------------               
    //  Clock Attributes
    //----------------------------------------------------------------------------------------------    
    .RXRECCLKOUT0_SEL                   ( 2'b00),
    .RXRECCLKOUT1_SEL                   ( 2'b00),                    

    //----------------------------------------------------------------------------------------------
    //  QPLL0 Attributes 
    //----------------------------------------------------------------------------------------------    
    .AEN_QPLL0_FBDIV                    (1'b1),                                 
    .QPLL0CLKOUT_RATE                   ("HALF"),                              
    .QPLL0_CFG0                         (16'b0011001100011100),                            
    .QPLL0_CFG1                         (16'b1101000000111000),                             
    .QPLL0_CFG1_G3                      (16'b1101000000111000),                             
    .QPLL0_CFG2                         (16'b0000111111000000),                             
    .QPLL0_CFG2_G3                      (16'b0000111111000000),                        
    .QPLL0_CFG3                         (16'b0000000100100000),                  
    .QPLL0_CFG4                         (16'b0000000011100111),
    .QPLL0_CP                           (10'b1111111111),                       // Optimized for PCIe PLL compliance
    .QPLL0_CP_G3                        (10'b0000011111),                       // Optimized for PCIe PLL compliance
    .QPLL0_FBDIV                        (QPLL_FBDIV),
    .QPLL0_FBDIV_G3                     (QPLL_FBDIV_G34),
    .QPLL0_INIT_CFG0                    (16'h02B2),
    .QPLL0_INIT_CFG1                    ( 8'b00000000),
    .QPLL0_LOCK_CFG                     (16'b0010010111101000),                             // [10] : 1'b1 = Auto VCO
    .QPLL0_LOCK_CFG_G3                  (16'b0010010111101000),                             // [10] : 1'b1 = Auto VCO
    .QPLL0_LPF                          (10'b0100110101),                       // Optimized for PCIe PLL compliance
    .QPLL0_LPF_G3                       (10'b1111111111),                       // Optimized for PCIe PLL compliance
    .QPLL0_PCI_EN                       ( 1'b1),                                
    .QPLL0_RATE_SW_USE_DRP              ( 1'b0),                                // Advance PCIe feature
    .QPLL0_REFCLK_DIV                   (1),
    .QPLL0_SDM_CFG0                     (16'b0000000011000000),                
    .QPLL0_SDM_CFG1                     (16'b0000000000000000),
    .QPLL0_SDM_CFG2                     (16'b0000000000000000),
                     
    //---------------------------------------------------------------------------------------------- 
    //  QPLL1 Attributes               
    //----------------------------------------------------------------------------------------------    
    .AEN_QPLL1_FBDIV                    (1'b1),                                 
    .QPLL1CLKOUT_RATE                   ("HALF"),                              
    .QPLL1_CFG0                         (16'b0011001100011100),                             
    .QPLL1_CFG1                         (16'b0001000000101000),                             
    .QPLL1_CFG1_G3                      (16'b0001000000101000),                             
    .QPLL1_CFG2                         (16'b0000111111000011),                             
    .QPLL1_CFG2_G3                      (16'b0000000100100000),                         
    .QPLL1_CFG3                         (16'b0000000100100000),                  
    .QPLL1_CFG4                         (16'b0000000001100011),
    .QPLL1_CP                           (10'b0100010101),                       // Optimized for PCIe PLL compliance
    .QPLL1_CP_G3                        (10'b0100010101),                       // Optimized for PCIe PLL compliance
    .QPLL1_FBDIV                        (QPLL_FBDIV),
    .QPLL1_FBDIV_G3                     (QPLL_FBDIV_G34),
    .QPLL1_INIT_CFG0                    (16'h02B2),
    .QPLL1_INIT_CFG1                    ( 8'b00000000),
    .QPLL1_LOCK_CFG                     (16'b0010010111101000),                             // [10] : 1'b1 = Auto VCO
    .QPLL1_LOCK_CFG_G3                  (16'b0010010111101000),                             // [10] : 1'b1 = Auto VCO
    .QPLL1_LPF                          (10'b0000010101),                       // Optimized for PCIe PLL compliance
    .QPLL1_LPF_G3                       (10'b0000010101),                       // Optimized for PCIe PLL compliance
    .QPLL1_PCI_EN                       ( 1'b1),                               
    .QPLL1_RATE_SW_USE_DRP              ( 1'b0),                                // Advance PCIe feature
    .QPLL1_REFCLK_DIV                   (1),
    .QPLL1_SDM_CFG0                     (16'b0000000011000000),                 
    .QPLL1_SDM_CFG1                     (16'b0000000000000000),
    .QPLL1_SDM_CFG2                     (16'b0000000000000000),
 
    //----------------------------------------------------------------------------------------------
    //  PPF Attributes                                                         
    //----------------------------------------------------------------------------------------------      
    .PPF0_CFG                           (16'h0FFF),                            
    .PPF1_CFG                           (16'h0FFF),                           
    
    //----------------------------------------------------------------------------------------------
    //  Bias Attributes                                                          
    //----------------------------------------------------------------------------------------------
    .BIAS_CFG0                          (16'b0000000000000000),
    .BIAS_CFG1                          (16'b0000000000000000),
    .BIAS_CFG2                          (16'b0000000100100100),                 // Optimized for PCIe PLL compliance
    .BIAS_CFG3                          (16'b0000000001000001),                 
    .BIAS_CFG4                          (16'b0000000000010000),    
    .BIAS_CFG_RSVD                      (10'b0000000000),  
       
    //---------------------------------------------------------------------------------------------- 
    //  SDM0 Attributes                                                          
    //----------------------------------------------------------------------------------------------
    .A_SDM0TOGGLE                       ( 1'b0),
    .AEN_SDM0TOGGLE                     ( 1'b0),
    .SDM0INITSEED0_0                    (16'b0000000000000000),
    .SDM0INITSEED0_1                    ( 9'b000000000),
    
    //---------------------------------------------------------------------------------------------- 
    //  SDM1 Attributes                                                          
    //----------------------------------------------------------------------------------------------     
    .A_SDM1DATA_HIGH                    ( 9'b000000000),
    .A_SDM1DATA_LOW                     (16'b0000000000000000),
    .A_SDM1TOGGLE                       ( 1'b0),
    .AEN_SDM1TOGGLE                     ( 1'b0),
    .SDM1INITSEED0_0                    (16'b0000000000000000),
    .SDM1INITSEED0_1                    ( 9'b000000000),     
          
    //----------------------------------------------------------------------------------------------
    //  Reserved & MISC Attributes                                                         
    //----------------------------------------------------------------------------------------------            
    .COMMON_CFG0                        (16'b0000000000000000),
    .COMMON_CFG1                        (16'b0000000000000000),
    .POR_CFG                            (16'b0000000000000000),                 // CHECK      
    .RSVD_ATTR0                         (16'b0000000000000000),                 // CHECK
    .RSVD_ATTR1                         (16'b0000000000000000),    
    .RSVD_ATTR2                         (16'b0000000000000000),                 // CHECK                
    .RSVD_ATTR3                         (16'b0000000000000000),
    .SARC_ENB                           ( 1'b0),
    .SARC_SEL                           ( 1'b0)
)
gthe4_common_smsw_i 
(       
    //----------------------------------------------------------------------------------------------
    //  QPLL0 Clock Ports
    //----------------------------------------------------------------------------------------------
    .GTGREFCLK0                         ( 1'd0), 
    .GTREFCLK00                         (GTCOM_REFCLK),                         
    .GTREFCLK10                         ( 1'd0),
    .GTNORTHREFCLK00                    ( 1'd0),
    .GTNORTHREFCLK10                    ( 1'd0),
    .GTSOUTHREFCLK00                    ( 1'd0),
    .GTSOUTHREFCLK10                    ( 1'd0),
   
    .REFCLKOUTMONITOR0                  (),
    .RXRECCLK0SEL                       (),
    
    //----------------------------------------------------------------------------------------------
    //  QPLL1 Clock Ports
    //----------------------------------------------------------------------------------------------
    .GTGREFCLK1                         ( 1'd0),
    .GTREFCLK01                         (GTCOM_REFCLK),
    .GTREFCLK11                         ( 1'd0),
    .GTNORTHREFCLK01                    ( 1'd0),    
    .GTNORTHREFCLK11                    ( 1'd0),
    .GTSOUTHREFCLK01                    ( 1'd0),
    .GTSOUTHREFCLK11                    ( 1'd0),        
        
    .REFCLKOUTMONITOR1                  (),  
    .RXRECCLK1SEL	                      (), 
        
    //----------------------------------------------------------------------------------------------
    //  QPLL0 Ports
    //----------------------------------------------------------------------------------------------
    .QPLL0CLKRSVD0                      ( 1'd0),
    .QPLL0CLKRSVD1                      ( 1'd0),                              
    .QPLL0FBDIV                         ( 8'd0),                                // CHECK
    .QPLL0LOCKDETCLK                    ( 1'd0),
    .QPLL0LOCKEN                        ( 1'd1),
    .QPLL0PD                            (GTCOM_QPLL0PD),                        
    .QPLL0REFCLKSEL                     ( 3'd1),                                                          
    .QPLL0RESET                         (GTCOM_QPLL0RESET),                     
       
    .QPLL0FBCLKLOST                     (),
    .QPLL0LOCK                          (GTCOM_QPLL0LOCK),
    .QPLL0OUTCLK                        (GTCOM_QPLL0OUTCLK),
    .QPLL0OUTREFCLK                     (GTCOM_QPLL0OUTREFCLK),
    .QPLL0REFCLKLOST                    (),     
    .QPLLDMONITOR0                      (),                                                                      
                                               
    //----------------------------------------------------------------------------------------------
    //  QPLL1 Ports
    //----------------------------------------------------------------------------------------------
    .QPLL1CLKRSVD0                      ( 1'd0),
    .QPLL1CLKRSVD1                      ( 1'd0),                                
    .QPLL1FBDIV                         ( 8'd0),                                // CHECK
    .QPLL1LOCKDETCLK                    ( 1'd0),
    .QPLL1LOCKEN                        ( 1'd1),
    .QPLL1PD                            (GTCOM_QPLL1PD),
    .QPLL1REFCLKSEL                     ( 3'd1),                        
    .QPLL1RESET                         (GTCOM_QPLL1RESET),      
     
    .QPLL1FBCLKLOST                     (),  
    .QPLL1LOCK                          (GTCOM_QPLL1LOCK),       
    .QPLL1OUTCLK                        (GTCOM_QPLL1OUTCLK),     
    .QPLL1OUTREFCLK                     (GTCOM_QPLL1OUTREFCLK),                       
    .QPLL1REFCLKLOST                    (),  
    .QPLLDMONITOR1                      (),            
         
    //----------------------------------------------------------------------------------------------
    //  PCIe Ports
    //----------------------------------------------------------------------------------------------
    .PCIERATEQPLL0                      (GTCOM_QPLLRATE),           
    .PCIERATEQPLL1                      (GTCOM_QPLLRATE),       
                                                                                                       
    //----------------------------------------------------------------------------------------------
    //  DRP Ports
    //----------------------------------------------------------------------------------------------
    .DRPCLK                             (GTCOM_DRPCLK),                                        
    .DRPADDR                            (GTCOM_DRPADDR),                                       
    .DRPEN                              (GTCOM_DRPEN),                                             
    .DRPWE                              (GTCOM_DRPWE),     
    .DRPDI                              (GTCOM_DRPDI),                                      
                                                                         
    .DRPRDY                             (GTCOM_DRPRDY),    
    .DRPDO                              (GTCOM_DRPDO),                                      
        
    //----------------------------------------------------------------------------------------------
    //  rCal Ports
    //----------------------------------------------------------------------------------------------        
    .RCALENB                            ( 1'd1),          
                                                                                                        
    //----------------------------------------------------------------------------------------------
    //  Band Gap Ports
    //----------------------------------------------------------------------------------------------
    .BGBYPASSB                          ( 1'b1),                                
    .BGMONITORENB                       ( 1'b1),                                
    .BGPDB                              ( 1'b1),  
    .BGRCALOVRD                         ( 5'b11111),                                 
    .BGRCALOVRDENB                      ( 1'b1),                                                            
        
    //----------------------------------------------------------------------------------------------
    //  SDM0 Ports
    //----------------------------------------------------------------------------------------------
    .SDM0DATA                           (25'd0),
    .SDM0RESET                          ( 1'd0),
    .SDM0TOGGLE                         ( 1'd0), 
    .SDM0WIDTH                          ( 2'd0),
    
    .SDM0FINALOUT                       (),
    .SDM0TESTDATA                       (),

    //----------------------------------------------------------------------------------------------
    //  SDM1 Ports
    //----------------------------------------------------------------------------------------------
    .SDM1DATA                           (25'd0),
    .SDM1RESET                          ( 1'd0),
    .SDM1TOGGLE                         ( 1'd0), 
    .SDM1WIDTH                          ( 2'd0),
    
    .SDM1FINALOUT                       (),
    .SDM1TESTDATA                       (),

    //----------------------------------------------------------------------------------------------
    //  TCON Ports
    //----------------------------------------------------------------------------------------------
    .TCONGPI                            (10'd0),
    .TCONPOWERUP                        ( 1'd0),
    .TCONRESET                          ( 2'd0),
    .TCONRSVDIN1                        ( 2'd0),
    
    .TCONGPO                            (),
    .TCONRSVDOUT0                       (),

    //----------------------------------------------------------------------------------------------
    //  Reserved & MISC Ports
    //----------------------------------------------------------------------------------------------
    .PMARSVD0                           ( 8'd0),            
    .PMARSVD1                           ( 8'd0),  
    .QPLLRSVD1                          ( 8'd0),
    .QPLLRSVD2                          ( 5'd0),               
    .QPLLRSVD3                          ( 5'd0),          
    .QPLLRSVD4                          ( 8'd0),                   

    .PMARSVDOUT0                        (),
    .PMARSVDOUT1                        ()
);
end
endgenerate

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_gt_phy_clk.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
//  Design :  PHY Wrapper 
//  Module :  PHY Clock
//--------------------------------------------------------------------------------------------------

`timescale 1ps / 1ps

//--------------------------------------------------------------------------------------------------
//  PHY Clock Module
//--------------------------------------------------------------------------------------------------
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_gt_phy_clk #
(
    parameter integer PHY_MAX_SPEED     = 4, 
    parameter         PHY_GEN4_64BIT_EN = "FALSE",
    parameter integer PHY_CORECLK_FREQ  = 2,  
    parameter integer PHY_USERCLK_FREQ  = 4, 
    parameter integer PHY_MCAPCLK_FREQ  = 4          
)
(
    //--------------------------------------------------------------------------
    //  CLK Port
    //--------------------------------------------------------------------------
    input                               CLK_TXOUTCLK,
    output                              CLK_PCLK2_GT,

    //--------------------------------------------------------------------------
    //  PCLK Ports
    //--------------------------------------------------------------------------
    input                               CLK_PCLK_CE,
    input                               CLK_PCLK_CEMASK,
    input                               CLK_PCLK_CLR,
    input                               CLK_PCLK_CLRMASK,
    input       [ 2:0]                  CLK_PCLK_DIV,
    output                              CLK_PCLK,
    
    //--------------------------------------------------------------------------
    //  PCLK2 Ports
    //--------------------------------------------------------------------------
    input                               CLK_PCLK2_CE,
    input                               CLK_PCLK2_CEMASK,
    input                               CLK_PCLK2_CLR,
    input                               CLK_PCLK2_CLRMASK,
    input       [ 2:0]                  CLK_PCLK2_DIV,
    output                              CLK_PCLK2,
    
    //--------------------------------------------------------------------------
    //  CORECLK Ports
    //--------------------------------------------------------------------------
    input                               CLK_CORECLK_CE,
    input                               CLK_CORECLK_CEMASK,
    input                               CLK_CORECLK_CLR,
    input                               CLK_CORECLK_CLRMASK,
    output                              CLK_CORECLK,      
    
    //--------------------------------------------------------------------------
    //  USERCLK Ports
    //--------------------------------------------------------------------------
    input                               CLK_USERCLK_CE,
    input                               CLK_USERCLK_CEMASK,
    input                               CLK_USERCLK_CLR,
    input                               CLK_USERCLK_CLRMASK,
    output                              CLK_USERCLK,    
    
    //--------------------------------------------------------------------------
    //  MCAPCLK Ports
    //--------------------------------------------------------------------------
    input                               CLK_MCAPCLK_CE,
    input                               CLK_MCAPCLK_CEMASK,
    input                               CLK_MCAPCLK_CLR,
    input                               CLK_MCAPCLK_CLRMASK,
    output                              CLK_MCAPCLK    
);
    //--------------------------------------------------------------------------
    //  Internal Signals
    //--------------------------------------------------------------------------                                     
    wire                                pclk;                                                                 
    wire                                pclk2;



    //----------------------------------------------------------------------------------------------
    //  Divider for CORECLK
    //----------------------------------------------------------------------------------------------     
    localparam [ 2:0] CORECLK_DIV_250MHZ = 3'd0;                                                    // 250.0 MHz
    localparam [ 2:0] CORECLK_DIV_500MHZ = (PHY_CORECLK_FREQ == 1) ? 3'd1 : 3'd0;                   // 250.0 MHZ : Default = 500.0 MHz                                
    
    localparam [ 2:0] CORECLK_DIV        = (PHY_MAX_SPEED     < 3) ? CORECLK_DIV_250MHZ : 
                                           (PHY_MAX_SPEED    == 4) ? CORECLK_DIV_500MHZ : 
                                           (PHY_CORECLK_FREQ == 1) ? CORECLK_DIV_250MHZ : CORECLK_DIV_500MHZ;



    //----------------------------------------------------------------------------------------------
    //  Divider for USERCLK
    //---------------------------------------------------------------------------------------------- 
    localparam [ 2:0] USERCLK_DIV_250MHZ = (PHY_USERCLK_FREQ == 3) ? 3'd0 :                         // 250.0 MHz
                                           (PHY_USERCLK_FREQ == 2) ? 3'd1 :                         // 125.0 MHz
                                           (PHY_USERCLK_FREQ == 1) ? 3'd3 : 3'd0;                   //  62.5 MHz : Default = 250.0 MHz
   
    localparam [ 2:0] USERCLK_DIV_500MHZ = (PHY_USERCLK_FREQ == 4) ? 3'd0 :                         // 500.0 MHz
                                           (PHY_USERCLK_FREQ == 3) ? 3'd1 :                         // 250.0 MHz
                                           (PHY_USERCLK_FREQ == 2) ? 3'd3 :                         // 125.0 MHz
                                           (PHY_USERCLK_FREQ == 1) ? 3'd7 : 3'd0;                   //  62.5 MHz : Default = 500.0 MHz
    
    localparam [ 2:0] USERCLK_DIV        = (PHY_MAX_SPEED     < 3) ? USERCLK_DIV_250MHZ :
                                           (PHY_MAX_SPEED    == 4) ? USERCLK_DIV_500MHZ : 
                                           (PHY_CORECLK_FREQ == 1) ? USERCLK_DIV_250MHZ : USERCLK_DIV_500MHZ;


                                           
    //----------------------------------------------------------------------------------------------
    //  Divider for MCAPCLK
    //---------------------------------------------------------------------------------------------- 
    localparam [ 2:0] MCAPCLK_DIV_250MHZ = (PHY_MCAPCLK_FREQ == 3) ? 3'd0 :                         // 250.0 MHz
                                           (PHY_MCAPCLK_FREQ == 2) ? 3'd1 :                         // 125.0 MHz
                                           (PHY_MCAPCLK_FREQ == 1) ? 3'd3 : 3'd0;                   //  62.5 MHz : Default = 250.0 MHz
   
    localparam [ 2:0] MCAPCLK_DIV_500MHZ = (PHY_MCAPCLK_FREQ == 4) ? 3'd0 :                         // 500.0 MHz
                                           (PHY_MCAPCLK_FREQ == 3) ? 3'd1 :                         // 250.0 MHz
                                           (PHY_MCAPCLK_FREQ == 2) ? 3'd3 :                         // 125.0 MHz
                                           (PHY_MCAPCLK_FREQ == 1) ? 3'd7 : 3'd0;                   //  62.5 MHz : Default = 500.0 MHz
    
    localparam [ 2:0] MCAPCLK_DIV        = (PHY_MAX_SPEED     < 3) ? MCAPCLK_DIV_250MHZ :
                                           (PHY_MAX_SPEED    == 4) ? MCAPCLK_DIV_500MHZ : 
                                           (PHY_CORECLK_FREQ == 1) ? MCAPCLK_DIV_250MHZ : MCAPCLK_DIV_500MHZ;

                                           

//--------------------------------------------------------------------------------------------------
//  BUFG_GT for PCLK
//--------------------------------------------------------------------------------------------------
BUFG_GT bufg_gt_pclk 
(
     //-------------------------------------------------------------------------
     //  Input Ports
     //-------------------------------------------------------------------------
    .CE                                 (CLK_PCLK_CE),
    .CEMASK                             (CLK_PCLK_CEMASK),
    .CLR                                (CLK_PCLK_CLR),
    .CLRMASK                            (CLK_PCLK_CLRMASK),
    .DIV                                (CLK_PCLK_DIV),
    .I                                  (CLK_TXOUTCLK),
    
     //-------------------------------------------------------------------------
     //  Output Ports
     //-------------------------------------------------------------------------
    .O                                  (pclk)
);



 assign pclk2 = pclk;


//--------------------------------------------------------------------------------------------------
//  BUFG_GT for CORECLK
//--------------------------------------------------------------------------------------------------
BUFG_GT bufg_gt_coreclk 
(
     //-------------------------------------------------------------------------
     //  Input Ports
     //-------------------------------------------------------------------------
    .CE                                 (CLK_CORECLK_CE),
    .CEMASK                             (CLK_CORECLK_CEMASK),
    .CLR                                (CLK_CORECLK_CLR),
    .CLRMASK                            (CLK_CORECLK_CLRMASK),
    .DIV                                (    CORECLK_DIV),
    .I                                  (CLK_TXOUTCLK),

     //-------------------------------------------------------------------------
     //  Output Ports
     //-------------------------------------------------------------------------
    .O                                  (CLK_CORECLK)
);



//--------------------------------------------------------------------------------------------------
//  BUFG_GT for USERCLK
//--------------------------------------------------------------------------------------------------
BUFG_GT bufg_gt_userclk 
(
     //-------------------------------------------------------------------------
     //  Input Ports
     //-------------------------------------------------------------------------
    .CE                                 (CLK_USERCLK_CE),
    .CEMASK                             (CLK_USERCLK_CEMASK),
    .CLR                                (CLK_USERCLK_CLR),
    .CLRMASK                            (CLK_USERCLK_CLRMASK),
    .DIV                                (    USERCLK_DIV),
    .I                                  (CLK_TXOUTCLK),
    
     //-------------------------------------------------------------------------
     //  Output Ports
     //-------------------------------------------------------------------------
    .O                                  (CLK_USERCLK)
);



//--------------------------------------------------------------------------------------------------
//  BUFG_GT for MCAPCLK
//--------------------------------------------------------------------------------------------------
BUFG_GT bufg_gt_mcapclk
(
     //-------------------------------------------------------------------------
     //  Input Ports
     //-------------------------------------------------------------------------
    .CE                                 (CLK_MCAPCLK_CE),
    .CEMASK                             (CLK_MCAPCLK_CEMASK),
    .CLR                                (CLK_MCAPCLK_CLR),
    .CLRMASK                            (CLK_MCAPCLK_CLRMASK),
    .DIV                                (    MCAPCLK_DIV),
    .I                                  (CLK_TXOUTCLK),

     //-------------------------------------------------------------------------
     //  Output Ports
     //-------------------------------------------------------------------------
    .O                                  (CLK_MCAPCLK)
);


//--------------------------------------------------------------------------------------------------
//  PHY Clock Output
//--------------------------------------------------------------------------------------------------
assign CLK_PCLK     = pclk;
assign CLK_PCLK2    = pclk2;
assign CLK_PCLK2_GT = (PHY_GEN4_64BIT_EN == "TRUE") ? pclk2 : pclk;



endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_gt_phy_rst.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
//  Design :  PHY Wrapper
//  Module :  PHY Reset 
//--------------------------------------------------------------------------------------------------

`timescale 1ps / 1ps

//--------------------------------------------------------------------------------------------------
//  PHY Reset Module
//--------------------------------------------------------------------------------------------------
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_gt_phy_rst #
(
    parameter integer PHY_LANE      = 16,   
    parameter integer PHY_MAX_SPEED = 4,
    parameter integer SYNC_STAGE    = 3
)
(
    //-------------------------------------------------------------------------- 
    //  Input Ports
    //-------------------------------------------------------------------------- 
    input                               RST_REFCLK,
    input                               RST_PCLK,
    input                               RST_N,
    input       [PHY_LANE-1:0]          RST_GTPOWERGOOD,
    input       [PHY_LANE-1:0]          RST_CPLLLOCK,
    input       [(PHY_LANE-1)>>2:0]     RST_QPLL0LOCK,   
    input       [(PHY_LANE-1)>>2:0]     RST_QPLL1LOCK,
    input       [PHY_LANE-1:0]          RST_TXPROGDIVRESETDONE,
    input       [PHY_LANE-1:0]          RST_TXRESETDONE,    
    input       [PHY_LANE-1:0]          RST_RXRESETDONE, 
    input       [PHY_LANE-1:0]          RST_TXSYNC_DONE,   
    input       [PHY_LANE-1:0]          RST_PHYSTATUS,
    
    //-------------------------------------------------------------------------- 
    //  Output Ports
    //-------------------------------------------------------------------------- 
    output                              RST_RRST_N,
    output                              RST_PRST_N,
    output                              RST_CPLLPD,
    output                              RST_CPLLRESET,
    output                              RST_QPLLPD,
    output                              RST_QPLLRESET,
    output                              RST_TXPROGDIVRESET,
    output                              RST_GTRESET,
    output                              RST_USERRDY,
    output                              RST_TXSYNC_START,
    output                              RST_IDLE
);
    //-------------------------------------------------------------------------- 
    //  Reset Synchronized Signals
    //-------------------------------------------------------------------------- 
    (* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *) reg [ 3:0] rrst_n_r;
    (* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *) reg [ 3:0] prst_n_r;

    wire                                rrst_n;                                     
    wire                                prst_n;  
       
    //--------------------------------------------------------------------------
    //  Synchronized Signals
    //--------------------------------------------------------------------------                                     
    wire        [PHY_LANE-1:0]          gtpowergood_r;                                                                 
    wire        [PHY_LANE-1:0]          cplllock_r;
    wire        [(PHY_LANE-1)>>2:0]     qpll0lock_r;
    wire        [(PHY_LANE-1)>>2:0]     qpll1lock_r;
    wire        [PHY_LANE-1:0]          txprogdivresetdone_r;
    wire        [PHY_LANE-1:0]          txresetdone_r;  
    wire        [PHY_LANE-1:0]          rxresetdone_r;
    wire        [PHY_LANE-1:0]          txsync_done_r;
    wire        [PHY_LANE-1:0]          phystatus_r;
    
    //--------------------------------------------------------------------------
    //  Internal Signals
    //--------------------------------------------------------------------------
    wire                                gtpowergood_a;
    wire                                cplllock_a;
    wire                                qplllock_a;
    wire                                txprogdivresetdone_a;
    wire                                resetdone_a;
    wire                                txsync_done_a;
    wire                                phystatus_a;
    
    reg         [ 1:0]                  txsync_start_cnt;
    
    //--------------------------------------------------------------------------
    //  Output Delayed Signals
    //--------------------------------------------------------------------------     
    reg         [ 3:0]                  cpllpd_r;
    reg         [ 3:0]                  cpllreset_r;                                  
    reg         [ 3:0]                  qpllpd_r;
    reg         [ 3:0]                  qpllreset_r;                                
    reg         [ 3:0]                  txprogdivreset_r;
    reg         [ 3:0]                  gtreset_r;
    reg         [ 3:0]                  userrdy_r;
                
    wire                                cpllpd_dly;
    wire                                cpllreset_dly;                                    
    wire                                qpllpd_dly;
    wire                                qpllreset_dly;                        
    wire                                txprogdivreset_dly;
    wire                                gtreset_dly;
    wire                                userrdy_dly;
     
    //-------------------------------------------------------------------------- 
    //  FSM Signals
    //-------------------------------------------------------------------------- 
    reg [ 2:0] fsm;
    
    reg                                 idle;     
    reg                                 cpllpd;
    reg                                 cpllreset;
    reg                                 qpllpd;
    reg                                 qpllreset;
    reg                                 txprogdivreset;
    reg                                 gtreset;
    reg                                 userrdy; 
    reg                                 txsync_start;         
   
    //--------------------------------------------------------------------------
    //  FSM Encoding
    //-------------------------------------------------------------------------- 
    localparam FSM_IDLE               = 3'd0;
    localparam FSM_GTPOWERGOOD        = 3'd1;
    localparam FSM_PLLLOCK            = 3'd2;
    localparam FSM_TXPROGDIVRESETDONE = 3'd3;
    localparam FSM_RESETDONE          = 3'd4;
    localparam FSM_TXSYNC_START       = 3'd5;
    localparam FSM_TXSYNC_DONE        = 3'd6;
    localparam FSM_PHYSTATUS          = 3'd7;



//--------------------------------------------------------------------------------------------------
//  Reset Synchronizer for REFCLK
//--------------------------------------------------------------------------------------------------
always @ (posedge RST_REFCLK or negedge RST_N)
begin

    if (!RST_N) 
        rrst_n_r <= 4'd0;
    else
        rrst_n_r <= {rrst_n_r[2:0], 1'd1}; 
          
end   
 
assign rrst_n = rrst_n_r[3];



//--------------------------------------------------------------------------------------------------
//  Reset Synchronizer for PCLK
//--------------------------------------------------------------------------------------------------
always @ (posedge RST_PCLK or negedge RST_N)
begin

    if (!RST_N) 
        prst_n_r <= 4'd0;
    else
        prst_n_r <= {prst_n_r[2:0], 1'd1};
          
end   

assign prst_n = prst_n_r[3];



//--------------------------------------------------------------------------------------------------
//  Input Synchronizer or Pipeline
//--------------------------------------------------------------------------------------------------
xp4_usp_smsw_sync #(.WIDTH (PHY_LANE),            .STAGE (SYNC_STAGE)) sync_gtpowergood        (.CLK (RST_REFCLK), .D (RST_GTPOWERGOOD),        .Q (gtpowergood_r));
xp4_usp_smsw_sync #(.WIDTH (PHY_LANE),            .STAGE (SYNC_STAGE)) sync_cplllock           (.CLK (RST_REFCLK), .D (RST_CPLLLOCK),           .Q (cplllock_r));
xp4_usp_smsw_sync #(.WIDTH (((PHY_LANE-1)>>2)+1), .STAGE (SYNC_STAGE)) sync_qpll0lock          (.CLK (RST_REFCLK), .D (RST_QPLL0LOCK),          .Q (qpll0lock_r));
xp4_usp_smsw_sync #(.WIDTH (((PHY_LANE-1)>>2)+1), .STAGE (SYNC_STAGE)) sync_qpll1lock          (.CLK (RST_REFCLK), .D (RST_QPLL1LOCK),          .Q (qpll1lock_r));
xp4_usp_smsw_sync #(.WIDTH (PHY_LANE),            .STAGE (SYNC_STAGE)) sync_txprogdivresetdone (.CLK (RST_REFCLK), .D (RST_TXPROGDIVRESETDONE), .Q (txprogdivresetdone_r));
xp4_usp_smsw_sync #(.WIDTH (PHY_LANE),            .STAGE (SYNC_STAGE)) sync_txresetdone        (.CLK (RST_REFCLK), .D (RST_TXRESETDONE),        .Q (txresetdone_r));  
xp4_usp_smsw_sync #(.WIDTH (PHY_LANE),            .STAGE (SYNC_STAGE)) sync_rxresetdone        (.CLK (RST_REFCLK), .D (RST_RXRESETDONE),        .Q (rxresetdone_r));
xp4_usp_smsw_sync #(.WIDTH (PHY_LANE),            .STAGE (SYNC_STAGE)) sync_txsync_done        (.CLK (RST_REFCLK), .D (RST_TXSYNC_DONE),        .Q (txsync_done_r)); 
xp4_usp_smsw_sync #(.WIDTH (PHY_LANE),            .STAGE (SYNC_STAGE)) sync_phystatus          (.CLK (RST_REFCLK), .D (RST_PHYSTATUS),          .Q (phystatus_r));



//--------------------------------------------------------------------------------------------------
//  Convert per-lane signals to per-design 
//--------------------------------------------------------------------------------------------------
assign gtpowergood_a        = &gtpowergood_r;
assign cplllock_a           = (PHY_MAX_SPEED  < 3) ? (&cplllock_r)  : cplllock_r[0];
assign qplllock_a           = (PHY_MAX_SPEED == 4) ? (&qpll0lock_r) : (&qpll1lock_r);
assign txprogdivresetdone_a = &txprogdivresetdone_r;
assign resetdone_a          = (&txresetdone_r) && (&rxresetdone_r);
assign txsync_done_a        = &txsync_done_r;
assign phystatus_a          = |phystatus_r;                 



//--------------------------------------------------------------------------------------------------
//  TX Sync Alignment Start Counter
//--------------------------------------------------------------------------------------------------
always @ (posedge RST_REFCLK)
begin

    if (!rrst_n)
        txsync_start_cnt <= 2'd0;
    else
        if (fsm == FSM_TXSYNC_START)
            txsync_start_cnt <= txsync_start_cnt + 2'd1; 
        else
            txsync_start_cnt <= 2'd0;
            
end



//--------------------------------------------------------------------------------------------------
//  Reset FSM
//--------------------------------------------------------------------------------------------------
always @ (posedge RST_REFCLK)
begin

    if (!rrst_n)
        begin
        fsm            <= FSM_GTPOWERGOOD;
        idle           <= 1'd0;
        cpllpd         <= 1'd1;                               
        cpllreset      <= 1'd1;
        qpllpd         <= 1'd1;
        qpllreset      <= 1'd1;
        txprogdivreset <= 1'd1;
        gtreset        <= 1'd1;
        userrdy        <= 1'd0;
        txsync_start   <= 1'd0;
        end
    else
        begin
        
        case (fsm)
            
        //------------------------------------------------------------------------------------------
        //  Stay in IDLE state until system reset is released
        //------------------------------------------------------------------------------------------
        FSM_IDLE :
        
            begin
            if (!rrst_n)
                begin
                fsm            <= FSM_GTPOWERGOOD;
                idle           <= 1'd0;
                cpllpd         <= 1'd1;
                cpllreset      <= 1'd1;
                qpllpd         <= 1'd1;
                qpllreset      <= 1'd1;
                txprogdivreset <= 1'd1;
                gtreset        <= 1'd1;
                userrdy        <= 1'd0;
                txsync_start   <= 1'd0;
                end
            else
                begin
                fsm            <= FSM_IDLE;
                idle           <= 1'd1;
                cpllpd         <= cpllpd;
                cpllreset      <= cpllreset;
                qpllpd         <= qpllpd;
                qpllreset      <= qpllreset;
                txprogdivreset <= txprogdivreset;
                gtreset        <= gtreset;
                userrdy        <= userrdy;
                txsync_start   <= txsync_start;
                end
            end   
            
        //------------------------------------------------------------------------------------------
        //  Release [CPLL/QPLL]PD and wait for GTPOWERGOOD to assert HIGH
        //------------------------------------------------------------------------------------------
        FSM_GTPOWERGOOD :
        
            begin
            fsm            <= (gtpowergood_a && (!cplllock_a) && (!qplllock_a || PHY_MAX_SPEED < 3)) ? FSM_PLLLOCK : FSM_GTPOWERGOOD;
            idle           <= idle;
            cpllpd         <= 1'd0;
            cpllreset      <= cpllreset;
            qpllpd         <= (PHY_MAX_SPEED < 3) ? 1'd1 : 1'd0;
            qpllreset      <= qpllreset;
            txprogdivreset <= txprogdivreset;
            gtreset        <= gtreset;
            userrdy        <= userrdy;
            txsync_start   <= txsync_start;
            end    
            
        //------------------------------------------------------------------------------------------
        //  Release [CPLL/QPLL]RESET and wait for [CPLL/QPLL]LOCK to assert HIGH
        //------------------------------------------------------------------------------------------
        FSM_PLLLOCK :
        
            begin
            fsm            <= (cplllock_a && (qplllock_a || PHY_MAX_SPEED < 3)) ? FSM_TXPROGDIVRESETDONE : FSM_PLLLOCK;
            idle           <= idle;
            cpllpd         <= cpllpd;
            cpllreset      <= 1'd0;
            qpllpd         <= qpllpd;
            qpllreset      <= (PHY_MAX_SPEED < 3) ? 1'd1 : 1'd0;
            txprogdivreset <= txprogdivreset;
            gtreset        <= gtreset;
            userrdy        <= userrdy;
            txsync_start   <= txsync_start;
            end

        //------------------------------------------------------------------------------------------
        //  Release TXPROGDIVRESET and wait for TXPROGDIVRESETDONE to assert HIGH
        //------------------------------------------------------------------------------------------
        FSM_TXPROGDIVRESETDONE :
        
            begin
            fsm            <= txprogdivresetdone_a ? FSM_RESETDONE : FSM_TXPROGDIVRESETDONE;  
            idle           <= idle;
            cpllpd         <= cpllpd;
            cpllreset      <= cpllreset;
            qpllpd         <= qpllpd;
            qpllreset      <= qpllreset;
            txprogdivreset <= 1'd0;
            gtreset        <= gtreset;
            userrdy        <= userrdy;
            txsync_start   <= txsync_start;
            end
            
        //------------------------------------------------------------------------------------------
        //  Release GT[TX/RX]RESET, assert [TX/RX]USERRDY, and wait for [TX/RX]RESETDONE to assert HIGH
        //------------------------------------------------------------------------------------------
        FSM_RESETDONE :
        
            begin
            fsm            <= resetdone_a ? FSM_TXSYNC_START : FSM_RESETDONE;  
            idle           <= idle;
            cpllpd         <= cpllpd;
            cpllreset      <= cpllreset;
            qpllpd         <= qpllpd;
            qpllreset      <= qpllreset;
            txprogdivreset <= txprogdivreset;
            gtreset        <= 1'd0;
            userrdy        <= 1'd1;
            txsync_start   <= txsync_start;
            end
        
        //------------------------------------------------------------------------------------------
        //  Start TX sync alignment.  Extend TXSYNC_START pulse by few REFCLK cycles
        //------------------------------------------------------------------------------------------
        FSM_TXSYNC_START :
        
            begin
            fsm            <= (!txsync_done_a && (txsync_start_cnt == 2'd3)) ? FSM_TXSYNC_DONE : FSM_TXSYNC_START;
            idle           <= idle;
            cpllpd         <= cpllpd;
            cpllreset      <= cpllreset;
            qpllpd         <= qpllpd;   
            qpllreset      <= qpllreset;
            txprogdivreset <= txprogdivreset;
            gtreset        <= gtreset;
            userrdy        <= userrdy;
            txsync_start   <= 1'd1;
            end
            
        //------------------------------------------------------------------------------------------
        //  Wait for TX sync alignment done
        //------------------------------------------------------------------------------------------
        FSM_TXSYNC_DONE :
        
            begin
            fsm            <= txsync_done_a ? FSM_PHYSTATUS : FSM_TXSYNC_DONE;
            idle           <= idle;
            cpllpd         <= cpllpd;
            cpllreset      <= cpllreset;
            qpllpd         <= qpllpd;
            qpllreset      <= qpllreset;
            txprogdivreset <= txprogdivreset;
            gtreset        <= gtreset;
            userrdy        <= userrdy;
            txsync_start   <= 1'd0;
            end    
            
        //------------------------------------------------------------------------------------------
        //  Wait for PHYSTATUS to de-assert LOW
        //------------------------------------------------------------------------------------------
        FSM_PHYSTATUS :
        
            begin
            fsm            <= !phystatus_a ? FSM_IDLE : FSM_PHYSTATUS;  
            idle           <= 1'd1;
            cpllpd         <= cpllpd;
            cpllreset      <= cpllreset;
            qpllpd         <= qpllpd;
            qpllreset      <= qpllreset;
            txprogdivreset <= txprogdivreset;
            gtreset        <= gtreset;
            userrdy        <= userrdy;
            txsync_start   <= txsync_start;
            end 
            
        //------------------------------------------------------------------------------------------
        //  Default State
        //------------------------------------------------------------------------------------------
        default :
        
            begin
            fsm            <= FSM_IDLE;
            idle           <= 1'd0;
            cpllpd         <= 1'd1;
            cpllreset      <= 1'd1;
            qpllpd         <= 1'd1;
            qpllreset      <= 1'd1;
            txprogdivreset <= 1'd1;
            gtreset        <= 1'd1;
            userrdy        <= 1'd0;
            txsync_start   <= 1'd0;
            end

        endcase
        
        end
        
end



//--------------------------------------------------------------------------------------------------
//  Delay Outputs
//--------------------------------------------------------------------------------------------------
always @ (posedge RST_REFCLK)
begin

    cpllpd_r         <= {cpllpd_r[2:0],         cpllpd}; 
    cpllreset_r      <= {cpllreset_r[2:0],      cpllreset}; 
    qpllpd_r         <= {qpllpd_r[2:0],         qpllpd}; 
    qpllreset_r      <= {qpllreset_r[2:0],      qpllreset}; 
    txprogdivreset_r <= {txprogdivreset_r[2:0], txprogdivreset}; 
    gtreset_r        <= {gtreset_r[2:0],        gtreset};    
    userrdy_r        <= {userrdy_r[2:0],        userrdy}; 
            
end

assign cpllpd_dly         = cpllpd_r[3];
assign cpllreset_dly      = cpllreset_r[3];
assign qpllpd_dly         = qpllpd_r[3];
assign qpllreset_dly      = qpllreset_r[3];
assign txprogdivreset_dly = txprogdivreset_r[3];
assign gtreset_dly        = gtreset_r[3];
assign userrdy_dly        = userrdy_r[3];



//--------------------------------------------------------------------------------------------------
//  PHY Reset Outputs
//--------------------------------------------------------------------------------------------------
assign RST_RRST_N         = rrst_n;
assign RST_PRST_N         = prst_n;

assign RST_CPLLPD         = cpllpd_dly;
assign RST_CPLLRESET      = cpllreset_dly; 
assign RST_QPLLPD         = qpllpd_dly;
assign RST_QPLLRESET      = qpllreset_dly;
assign RST_TXPROGDIVRESET = txprogdivreset_dly;
assign RST_GTRESET        = gtreset_dly;  
assign RST_USERRDY        = userrdy_dly;
assign RST_TXSYNC_START   = txsync_start;
assign RST_IDLE           = idle;



endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_gt_phy_rxeq.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
//  Design :  PHY Wrapper                                                             
//  Module :  RX Equalization                                                                   
//--------------------------------------------------------------------------------------------------

`timescale 1ps / 1ps
 
//--------------------------------------------------------------------------------------------------
//  RX Equalization Module
//--------------------------------------------------------------------------------------------------
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_gt_phy_rxeq #
(
    parameter         PHY_SIM_EN      = "FALSE",   
    parameter integer PHY_LP_TXPRESET = 4,
    parameter integer SYNC_STAGE      = 3                        
)
(
    //-------------------------------------------------------------------------- 
    //  Input Ports
    //-------------------------------------------------------------------------- 
    input                               RXEQ_CLK,                            
    input                               RXEQ_RST_N,
    
    input       [ 1:0]                  RXEQ_CTRL,    
    input       [ 2:0]                  RXEQ_PRESET,
    input       [ 3:0]                  RXEQ_TXPRESET,
    input       [ 5:0]                  RXEQ_TXCOEFF,
    input       [ 5:0]                  RXEQ_LFFS,
    
    //-------------------------------------------------------------------------- 
    //  Output Ports
    //-------------------------------------------------------------------------- 
    output                              RXEQ_LFFS_SEL, 
    output      [17:0]                  RXEQ_NEW_TXCOEFF,
    output                              RXEQ_ADAPT_DONE,
    output                              RXEQ_DONE 
);          
    //--------------------------------------------------------------------------
    //  Synchronized Signals
    //--------------------------------------------------------------------------   
    wire        [ 1:0]                  ctrl_r;
    wire        [ 2:0]                  preset_r;
    wire        [ 3:0]                  txpreset_r;
    wire        [ 5:0]                  txcoeff_r;
    wire        [ 5:0]                  lffs_r;

    //--------------------------------------------------------------------------
    //  Internal Signals
    //--------------------------------------------------------------------------
    reg         [ 21:0]                 adapt_cnt;

    //--------------------------------------------------------------------------
    //  FSM Signals                                                            
    //--------------------------------------------------------------------------    
    reg         [ 2:0]                  fsm;
    reg         [ 3:0]                  txpreset;
    reg         [17:0]                  txcoeff;
    reg         [ 1:0]                  txcoeff_cnt;
    reg                                 lffs_sel;
    reg                                 adapt_done;
    reg                                 adapt_2nd;
    reg                                 done;
   
    //----------------------------------------------------------------------------------------------  
    //  FSM Encoding                                                                                  
    //----------------------------------------------------------------------------------------------                                            
    localparam FSM_IDLE    = 3'd0; 
    localparam FSM_PRESET  = 3'd1;                                     
    localparam FSM_TXCOEFF = 3'd2;
    localparam FSM_ADAPT   = 3'd3;
    localparam FSM_DONE    = 3'd4;                                  

    //--------------------------------------------------------------------------
    //  New TX Coefficient
    //--------------------------------------------------------------------------
    localparam NEW_TXCOEFF = (PHY_LP_TXPRESET == 10) ? 18'd10 :
                             (PHY_LP_TXPRESET ==  9) ? 18'd9  :
                             (PHY_LP_TXPRESET ==  8) ? 18'd8  :
                             (PHY_LP_TXPRESET ==  7) ? 18'd7  :
                             (PHY_LP_TXPRESET ==  6) ? 18'd6  :                                                                     
                             (PHY_LP_TXPRESET ==  5) ? 18'd5  :
                             (PHY_LP_TXPRESET ==  4) ? 18'd4  :
                             (PHY_LP_TXPRESET ==  3) ? 18'd3  :
                             (PHY_LP_TXPRESET ==  2) ? 18'd2  :           
                             (PHY_LP_TXPRESET ==  1) ? 18'd1  :
                             (PHY_LP_TXPRESET ==  0) ? 18'd0  : 18'd0;   

    //--------------------------------------------------------------------------
    //  Counters (Simulation vs. Silicon)
    //--------------------------------------------------------------------------
    localparam ADAPT_MAX = (PHY_SIM_EN == "TRUE") ? 22'd1000 : 22'd2000000;
  
    
    
//--------------------------------------------------------------------------------------------------
//  Input Synchronizer
//--------------------------------------------------------------------------------------------------
xp4_usp_smsw_sync #(.WIDTH (2), .STAGE (SYNC_STAGE)) sync_ctrl     (.CLK (RXEQ_CLK), .D (RXEQ_CTRL),     .Q (ctrl_r));
xp4_usp_smsw_sync #(.WIDTH (3), .STAGE (SYNC_STAGE)) sync_preset   (.CLK (RXEQ_CLK), .D (RXEQ_PRESET),   .Q (preset_r));
xp4_usp_smsw_sync #(.WIDTH (4), .STAGE (SYNC_STAGE)) sync_txpreset (.CLK (RXEQ_CLK), .D (RXEQ_TXPRESET), .Q (txpreset_r));    
xp4_usp_smsw_sync #(.WIDTH (6), .STAGE (SYNC_STAGE)) sync_txcoeff  (.CLK (RXEQ_CLK), .D (RXEQ_TXCOEFF),  .Q (txcoeff_r));
xp4_usp_smsw_sync #(.WIDTH (6), .STAGE (SYNC_STAGE)) sync_lffs     (.CLK (RXEQ_CLK), .D (RXEQ_LFFS),     .Q (lffs_r));            



//--------------------------------------------------------------------------------------------------
//  Adaptation Counter
//--------------------------------------------------------------------------------------------------
always @ (posedge RXEQ_CLK)
begin

    if (!RXEQ_RST_N)
        begin
        adapt_cnt <= 22'd0;
        end
    else
        begin
        
        //----------------------------------------------------------------------
        //  Increment Counter
        //----------------------------------------------------------------------
        if (fsm == FSM_ADAPT)
            begin
            adapt_cnt <= adapt_cnt + 22'd1;
            end
            
        //----------------------------------------------------------------------
        //  Reset Counter
        //----------------------------------------------------------------------
        else
            begin
            adapt_cnt <= 22'd0;
            end

        end
        
end



//-------------------------------------------------------------------------------------------------- 
//  RX Equalization FSM                                                                              
//-------------------------------------------------------------------------------------------------- 
always @ (posedge RXEQ_CLK)
begin

    if (!RXEQ_RST_N)
        begin
        fsm         <= FSM_IDLE; 
        txpreset    <=  4'd0;
        txcoeff     <= 18'd0;
        txcoeff_cnt <=  2'd0;
        lffs_sel    <=  1'd0;
        adapt_done  <=  1'd0;
        adapt_2nd   <=  1'd1;
        done        <=  1'd0;
        end                    
    else
        begin
        
        case (fsm)
        
        //------------------------------------------------------------------------------------------
        //  Wait until RXEQ_CTRL != 2'b00
        //------------------------------------------------------------------------------------------
        FSM_IDLE :
        
            begin
            
            case (ctrl_r)
                
            //------------------------------------------------------------------
            //  Idle
            //------------------------------------------------------------------
            2'd0 :
            
                begin
                fsm         <= FSM_IDLE; 
                txpreset    <=  4'd0;
                txcoeff     <= 18'd0;
                txcoeff_cnt <=  2'd0;
                lffs_sel    <=  1'd0;
                adapt_done  <=  1'd0;
                adapt_2nd   <= adapt_2nd;
                done        <=  1'd0;
                end      
                
            //------------------------------------------------------------------
            //  Preset
            //------------------------------------------------------------------
            2'd1 :
            
                begin
                fsm         <= FSM_PRESET; 
                txpreset    <=  4'd0;
                txcoeff     <= 18'd0;
                txcoeff_cnt <=  2'd0;
                lffs_sel    <=  1'd0;
                adapt_done  <=  1'd0;
                adapt_2nd   <= adapt_2nd;
                done        <=  1'd0;
                end  
                
            //------------------------------------------------------------------
            //  Coeff : Latch C(-1) and TXPRESET
            //------------------------------------------------------------------
            2'd2 :
            
                begin
                fsm         <= FSM_TXCOEFF; 
                txpreset    <= txpreset_r;
                txcoeff     <= {txcoeff_r, txcoeff[17:6]};
                txcoeff_cnt <= 2'd1;
                lffs_sel    <= 1'd1;
                adapt_done  <= 1'd0;
                adapt_2nd   <= !adapt_2nd;                                      // Toggle adapt done
                done        <= 1'd0;
                end
                
            //------------------------------------------------------------------
            //  Bypass : Latch C(-1) and TXPRESET
            //------------------------------------------------------------------
            2'd3 :
            
                begin
                fsm         <= FSM_TXCOEFF; 
                txpreset    <= txpreset_r;
                txcoeff     <= {txcoeff_r, txcoeff[17:6]};
                txcoeff_cnt <= 2'd1;
                lffs_sel    <= 1'd1;
                adapt_done  <= 1'd0;
                adapt_2nd   <= 1'd1;
                done        <= 1'd0;
                end
                
            //------------------------------------------------------------------
            //  Default
            //------------------------------------------------------------------
            default :
            
                begin
                fsm         <= FSM_IDLE; 
                txpreset    <=  4'd0;
                txcoeff     <= 18'd0;
                txcoeff_cnt <=  2'd0;
                lffs_sel    <=  1'd0;
                adapt_done  <=  1'd0;
                adapt_2nd   <= adapt_2nd;
                done        <=  1'd0;
                end
                
            endcase
            
            end
            
        //------------------------------------------------------------------------------------------
        //  Go to DONE state (RXEQ preset not supported)
        //------------------------------------------------------------------------------------------
        FSM_PRESET :
        
            begin
            fsm         <= FSM_DONE;
            txpreset    <=  4'd0;
            txcoeff     <= 18'd0; 
            txcoeff_cnt <=  2'd0;
            lffs_sel    <=  1'd0;
            adapt_done  <=  1'd0;
            adapt_2nd   <= adapt_2nd;
            done        <=  1'd0; 
            end        
            
        //------------------------------------------------------------------------------------------
        //  Latch C(0) and C(+1)
        //------------------------------------------------------------------------------------------
        FSM_TXCOEFF :
        
            begin
            fsm         <= (txcoeff_cnt == 2'd2) ? FSM_ADAPT : FSM_TXCOEFF;
            txpreset    <= txpreset;
            txcoeff     <= {txcoeff_r, txcoeff[17:6]};
            txcoeff_cnt <= txcoeff_cnt + 2'd1;
            lffs_sel    <= 1'd0;
            adapt_done  <= 1'd0;
            adapt_2nd   <= adapt_2nd;
            done        <= 1'd0; 
            end
   
        //------------------------------------------------------------------------------------------
        //  Wait for adaptation timer 
        //------------------------------------------------------------------------------------------
        FSM_ADAPT :
        
            begin            
            fsm         <= (adapt_cnt == ADAPT_MAX) || (!adapt_2nd) ? FSM_DONE : FSM_ADAPT;
            txpreset    <= txpreset;
            txcoeff     <= txcoeff;
            txcoeff_cnt <= 2'd0;
            lffs_sel    <= 1'd0;
            adapt_done  <= 1'd0;
            adapt_2nd   <= adapt_2nd;
            done        <= 1'd0;
            end             
             
        //------------------------------------------------------------------------------------------
        //  Assert RXEQ_DONE until RXEQ_CTRL == 2'd0
        //------------------------------------------------------------------------------------------
        FSM_DONE :
        
            begin
            fsm         <= (ctrl_r == 2'd0) ? FSM_IDLE : FSM_DONE;
            txpreset    <= txpreset;
            txcoeff     <= txcoeff;
            txcoeff_cnt <= 2'd0;
            lffs_sel    <= ((ctrl_r == 2'd2) || (ctrl_r == 2'd3));
            adapt_done  <= ((ctrl_r == 2'd2) || (ctrl_r == 2'd3)) ? adapt_2nd : 1'd0;
            adapt_2nd   <= adapt_2nd;  
            done        <= 1'd1;
            end        
                          
        //------------------------------------------------------------------------------------------
        //  Default State
        //------------------------------------------------------------------------------------------
        default : 
        
            begin
            fsm         <= FSM_IDLE;
            txpreset    <=  4'd0;
            txcoeff     <= 18'd0;
            txcoeff_cnt <=  2'd0;
            lffs_sel    <=  1'd0;
            adapt_done  <=  1'd0; 
            adapt_2nd   <=  1'd1; 
            done        <=  1'd0; 
            end    
                    
        endcase
        
        end
        
end      



//-------------------------------------------------------------------------------------------------- 
//  RX Equalization Output                                                                           
//-------------------------------------------------------------------------------------------------- 
assign RXEQ_NEW_TXCOEFF = NEW_TXCOEFF;
assign RXEQ_LFFS_SEL    = lffs_sel;
assign RXEQ_ADAPT_DONE  = adapt_done;
assign RXEQ_DONE        = done;



endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_gt_phy_txeq.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
//  Design :  PCIe PHY Wrapper 
//  Module :  TX Equalization 
//--------------------------------------------------------------------------------------------------



`timescale 1ps / 1ps



//--------------------------------------------------------------------------------------------------
//  TX Equalization Module
//--------------------------------------------------------------------------------------------------
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_gt_phy_txeq #
(
    parameter integer PHY_GT_TXPRESET = 0,
    parameter integer SYNC_STAGE    = 3
)
(
    //-------------------------------------------------------------------------- 
    //  Input Ports
    //-------------------------------------------------------------------------- 
    input                               TXEQ_CLK,                            
    input                               TXEQ_RST_N,

    input       [ 1:0]                  TXEQ_CTRL,    
    input       [ 3:0]                  TXEQ_PRESET,
    input       [ 5:0]                  TXEQ_COEFF,
    
    //-------------------------------------------------------------------------- 
    //  Output Ports
    //-------------------------------------------------------------------------- 
    output  reg [ 4:0]                  TXEQ_PRECURSOR, 
    output  reg [ 6:0]                  TXEQ_MAINCURSOR,
    output  reg [ 4:0]                  TXEQ_POSTCURSOR,
    output  reg [17:0]                  TXEQ_NEW_COEFF,
    output  reg                         TXEQ_DONE
);          
    //--------------------------------------------------------------------------
    //  Synchronized Signals
    //-------------------------------------------------------------------------- 
    wire        [ 1:0]                  ctrl_r; 
    wire        [ 3:0]                  preset_r;
    wire        [ 5:0]                  coeff_r;
  
    //--------------------------------------------------------------------------
    //  Internal Signals
    //--------------------------------------------------------------------------
    reg         [18:0]                  preset;          
    reg                                 preset_done;
    
    //--------------------------------------------------------------------------
    //  FSM Signals                                                            
    //--------------------------------------------------------------------------    
    reg         [ 2:0]                  fsm;
    reg         [18:0]                  coeff;
    reg         [ 1:0]                  coeff_cnt;
    reg                                 done;
   
    //----------------------------------------------------------------------------------------------                   
    //  FSM Encoding                                                                               
    //----------------------------------------------------------------------------------------------                   
    localparam FSM_IDLE   = 3'd0; 
    localparam FSM_PRESET = 3'd1;                                     
    localparam FSM_COEFF  = 3'd2;
    localparam FSM_REMAP  = 3'd3;
    localparam FSM_QUERY  = 3'd4;                                     
    localparam FSM_DONE   = 3'd5;

    //----------------------------------------------------------------------------------------------
    //  TX Equalization Preset 
    //----------------------------------------------------------------------------------------------
    //  Advertise FS = 40
    //  Advertise LF = 12
    //  Actual    FS = 80
    //  Actual    LF = 24
    //----------------------------------------------------------------------------------------------
    //  Coefficient Rules:
    //  * C(-1) < Floor(FS/4)
    //  * C(-1) + C(0) + C(+1) = FS
    //  * C(0) - C(-1) - C(+1) >= LF
    //----------------------------------------------------------------------------------------------
    //  TXPRECURSOR  or C(-1) should be 20 or less
    //  TXMAINCURSOR or C( 0) should be 52 or more (automatically calcuated in GT)
    //  TXPOSTCURSOR or C(+1) should be 28 or less
    //----------------------------------------------------------------------------------------------                           
    localparam TXPRECURSOR_00  = 6'd0;   // 0.0 dB
    localparam TXMAINCURSOR_00 = 7'd58;                     
    localparam TXPOSTCURSOR_00 = 6'd22;  // 6.0 dB
                                         
    localparam TXPRECURSOR_01  = 6'd0;   // 0.0 dB
    localparam TXMAINCURSOR_01 = 7'd64;                               
    localparam TXPOSTCURSOR_01 = 6'd16;  // 3.5 dB
                                         
    localparam TXPRECURSOR_02  = 6'd0;   // 0.0 dB
    localparam TXMAINCURSOR_02 = 7'd62;                     
    localparam TXPOSTCURSOR_02 = 6'd18;  // 4.5 dB
                                         
    localparam TXPRECURSOR_03  = 6'd0;   // 0.0 dB
    localparam TXMAINCURSOR_03 = 7'd68;                     
    localparam TXPOSTCURSOR_03 = 6'd12;  // 2.5 dB
                                         
    localparam TXPRECURSOR_04  = 6'd0;   // 0.0 dB
    localparam TXMAINCURSOR_04 = 7'd80;                     
    localparam TXPOSTCURSOR_04 = 6'd0;   // 0.0 dB
                                         
    localparam TXPRECURSOR_05  = 6'd8;   // 2.0 dB
    localparam TXMAINCURSOR_05 = 7'd72;                     
    localparam TXPOSTCURSOR_05 = 6'd0;   // 0.0 dB
                                         
    localparam TXPRECURSOR_06  = 6'd10;  // 2.5 dB
    localparam TXMAINCURSOR_06 = 7'd70;                     
    localparam TXPOSTCURSOR_06 = 6'd0;   // 0.0 dB
                                         
    localparam TXPRECURSOR_07  = 6'd10;  // 3.5 dB
    localparam TXMAINCURSOR_07 = 7'd54;                     
    localparam TXPOSTCURSOR_07 = 6'd16;  // 6.0 dB
                                         
    localparam TXPRECURSOR_08  = 6'd12;  // 3.5 dB
    localparam TXMAINCURSOR_08 = 7'd56;                     
    localparam TXPOSTCURSOR_08 = 6'd12;  // 3.5 dB
                                         
    localparam TXPRECURSOR_09  = 6'd14;  // 3.5 dB
    localparam TXMAINCURSOR_09 = 7'd66;                    
    localparam TXPOSTCURSOR_09 = 6'd0;   // 0.0 dB
                                         
    localparam TXPRECURSOR_10  = 6'd0;   // 0.0 dB
    localparam TXMAINCURSOR_10 = 7'd54;                      
    localparam TXPOSTCURSOR_10 = 6'd26;  // 9.5 dB
    
//--------------------------------------------------------------------------------------------------
//  Input Synchronizer
//--------------------------------------------------------------------------------------------------
xp4_usp_smsw_sync #(.WIDTH (2), .STAGE (SYNC_STAGE)) sync_ctrl   (.CLK (TXEQ_CLK), .D (TXEQ_CTRL),   .Q (ctrl_r));
xp4_usp_smsw_sync #(.WIDTH (4), .STAGE (SYNC_STAGE)) sync_preset (.CLK (TXEQ_CLK), .D (TXEQ_PRESET), .Q (preset_r));
xp4_usp_smsw_sync #(.WIDTH (6), .STAGE (SYNC_STAGE)) sync_coeff  (.CLK (TXEQ_CLK), .D (TXEQ_COEFF),  .Q (coeff_r));



//--------------------------------------------------------------------------------------------------
//  TX Equalization Preset
//--------------------------------------------------------------------------------------------------
always @ (posedge TXEQ_CLK)
begin

    if (!TXEQ_RST_N)
        begin
        
        //------------------------------------------------------------------
        //  Default TX Equalization Preset                                 
        //------------------------------------------------------------------
        case (PHY_GT_TXPRESET)
            4'd0    : preset <= {TXPOSTCURSOR_00, TXMAINCURSOR_00, TXPRECURSOR_00};
            4'd1    : preset <= {TXPOSTCURSOR_01, TXMAINCURSOR_01, TXPRECURSOR_01};
            4'd2    : preset <= {TXPOSTCURSOR_02, TXMAINCURSOR_02, TXPRECURSOR_02};
            4'd3    : preset <= {TXPOSTCURSOR_03, TXMAINCURSOR_03, TXPRECURSOR_03};
            4'd4    : preset <= {TXPOSTCURSOR_04, TXMAINCURSOR_04, TXPRECURSOR_04};
            4'd5    : preset <= {TXPOSTCURSOR_05, TXMAINCURSOR_05, TXPRECURSOR_05};
            4'd6    : preset <= {TXPOSTCURSOR_06, TXMAINCURSOR_06, TXPRECURSOR_06};
            4'd7    : preset <= {TXPOSTCURSOR_07, TXMAINCURSOR_07, TXPRECURSOR_07};
            4'd8    : preset <= {TXPOSTCURSOR_08, TXMAINCURSOR_08, TXPRECURSOR_08};      
            4'd9    : preset <= {TXPOSTCURSOR_09, TXMAINCURSOR_09, TXPRECURSOR_09};   
            4'd10   : preset <= {TXPOSTCURSOR_10, TXMAINCURSOR_10, TXPRECURSOR_10};                 
            default : preset <= {TXPOSTCURSOR_00, TXMAINCURSOR_00, TXPRECURSOR_00};   
        endcase	       
        
        preset_done <= 1'd0;
        end                    
    else
        begin   
        if (fsm == FSM_PRESET)
            begin    
                
            //------------------------------------------------------------------
            //  Update TX Equalization Preset
            //------------------------------------------------------------------
            case (preset_r)
                4'd0    : preset <= {TXPOSTCURSOR_00, TXMAINCURSOR_00, TXPRECURSOR_00};
                4'd1    : preset <= {TXPOSTCURSOR_01, TXMAINCURSOR_01, TXPRECURSOR_01};
                4'd2    : preset <= {TXPOSTCURSOR_02, TXMAINCURSOR_02, TXPRECURSOR_02};
                4'd3    : preset <= {TXPOSTCURSOR_03, TXMAINCURSOR_03, TXPRECURSOR_03};
                4'd4    : preset <= {TXPOSTCURSOR_04, TXMAINCURSOR_04, TXPRECURSOR_04};
                4'd5    : preset <= {TXPOSTCURSOR_05, TXMAINCURSOR_05, TXPRECURSOR_05};
                4'd6    : preset <= {TXPOSTCURSOR_06, TXMAINCURSOR_06, TXPRECURSOR_06};
                4'd7    : preset <= {TXPOSTCURSOR_07, TXMAINCURSOR_07, TXPRECURSOR_07};
                4'd8    : preset <= {TXPOSTCURSOR_08, TXMAINCURSOR_08, TXPRECURSOR_08};      
                4'd9    : preset <= {TXPOSTCURSOR_09, TXMAINCURSOR_09, TXPRECURSOR_09}; 
                4'd10   : preset <= {TXPOSTCURSOR_10, TXMAINCURSOR_10, TXPRECURSOR_10};                   
                default : preset <= {TXPOSTCURSOR_00, TXMAINCURSOR_00, TXPRECURSOR_00};    
            endcase
              
            preset_done <= 1'd1;
            end
        else
            begin
            preset      <= preset;
            preset_done <= 1'd0;
            end
        end
        
end     



//--------------------------------------------------------------------------------------------------
//  TX Equalization FSM
//--------------------------------------------------------------------------------------------------
always @ (posedge TXEQ_CLK)
begin

    if (!TXEQ_RST_N)
        begin
        fsm       <= FSM_IDLE; 
        coeff     <= preset;
        coeff_cnt <= 2'd0;
        done      <= 1'd0;
        end                    
    else
        begin
        
        case (fsm)
        
        //------------------------------------------------------------------------------------------
        //  Wait until TXEQ_CTRL != 2'b00
        //------------------------------------------------------------------------------------------
        FSM_IDLE :
        
            begin
            done <= 1'd0;
            
            case (ctrl_r)
            
            //------------------------------------------------------------------
            //  Idle
            //------------------------------------------------------------------
            2'd0 :
            
                begin
                fsm       <= FSM_IDLE; 
                coeff     <= coeff;
                coeff_cnt <= 2'd0;
                end 
                
            //------------------------------------------------------------------
            //  Preset
            //------------------------------------------------------------------
            2'd1 :
            
                begin
                fsm       <= FSM_PRESET; 
                coeff     <= coeff;
                coeff_cnt <= 2'd0;
                end  
                
            //------------------------------------------------------------------
            //  Coeff : Latch C(-1) 
            //------------------------------------------------------------------
            2'd2 :
            
                begin
                fsm       <= FSM_COEFF; 
                coeff     <= {coeff_r, coeff[18:6]};
                coeff_cnt <= 2'd1;
                end
                
            //------------------------------------------------------------------
            //  Query
            //------------------------------------------------------------------
            2'd3 :
            
                begin
                fsm       <= FSM_QUERY; 
                coeff     <= coeff;
                coeff_cnt <= 2'd0;
                end
                
            //------------------------------------------------------------------
            //  Stay in IDLE state (Default)
            //------------------------------------------------------------------
            default :
            
                begin
                fsm       <= FSM_IDLE; 
                coeff     <= coeff;
                coeff_cnt <= 2'd0;
                end
                
            endcase
            
            end
            
        //------------------------------------------------------------------------------------------
        //  Wait for TXEQ preset done
        //------------------------------------------------------------------------------------------
        FSM_PRESET :
        
            begin
            fsm       <= preset_done ? FSM_DONE : FSM_PRESET;
            coeff     <= preset;
            coeff_cnt <= 2'd0;
            done      <= 1'd0;
            end    
            
        //------------------------------------------------------------------------------------------
        //  Latch C(0) and C(+1)
        //------------------------------------------------------------------------------------------
        FSM_COEFF :
        
            begin
            fsm <= (coeff_cnt == 2'd2) ? FSM_REMAP : FSM_COEFF;
            
            //------------------------------------------------------------------
            //  Shift in one extra bit for TXMAINCURSOR
            //------------------------------------------------------------------
            if (coeff_cnt == 2'd1)
                coeff <= {1'd0, coeff_r, coeff[18:7]};
            else
                coeff <= {coeff_r, coeff[18:6]};
                
            coeff_cnt <= coeff_cnt + 2'd1;
            done      <= 1'd0; 
            end
            
        //------------------------------------------------------------------------------------------
        //  Multiply coefficient by 2x
        //------------------------------------------------------------------------------------------
        FSM_REMAP :
        
            begin
            fsm       <= FSM_DONE;
            coeff     <= coeff << 1;        
            coeff_cnt <= 2'd0;
            done      <= 1'd0; 
            end
            
        //------------------------------------------------------------------------------------------
        //  Query to display current TXEQ_NEW_COEFF
        //------------------------------------------------------------------------------------------
        FSM_QUERY:
        
            begin
            fsm       <= FSM_DONE;
            coeff     <= coeff; 
            coeff_cnt <= 2'd0;
            done      <= 1'd0;
            end     
                  
        //------------------------------------------------------------------------------------------
        //  Assert TXEQ_DONE until TXEQ_CTRL == 2'd0
        //------------------------------------------------------------------------------------------
        FSM_DONE :
        
            begin
            fsm       <= (ctrl_r == 2'd0) ? FSM_IDLE : FSM_DONE;
            coeff     <= coeff;          
            coeff_cnt <= 2'd0;
            done      <= 1'd1;
            end        
                          
        //------------------------------------------------------------------------------------------
        //  Default State
        //------------------------------------------------------------------------------------------
        default : 
        
            begin
            fsm       <= FSM_IDLE;
            coeff     <= 19'd0; 
            coeff_cnt <=  2'd0;
            done      <=  1'd0;
            end    
                    
        endcase
        
        end
        
end  



//-------------------------------------------------------------------------------------------------- 
//  TX Equalization Output Register                                                                               
//-------------------------------------------------------------------------------------------------- 
always @ (posedge TXEQ_CLK)
begin

    if (!TXEQ_RST_N)
        begin
        TXEQ_PRECURSOR        <= coeff[ 4: 0];  
        TXEQ_MAINCURSOR       <= coeff[12: 6]; 
        TXEQ_POSTCURSOR       <= coeff[17:13];
        TXEQ_NEW_COEFF[17:12] <= {1'd0, coeff[18:14]};
        TXEQ_NEW_COEFF[11: 6] <= coeff[12:7]; 
        TXEQ_NEW_COEFF[ 5: 0] <= {1'd0, coeff[5:1]}; 
        TXEQ_DONE             <= 1'd0;
        end
    else           
        begin
        TXEQ_DONE <= done;
        
        //----------------------------------------------------------------------
        //  Divide TXEQ_NEW_COEFF by 2x and update output
        //----------------------------------------------------------------------
        if (fsm == FSM_DONE)
            begin
            TXEQ_PRECURSOR        <= coeff[ 4: 0]; 
            TXEQ_MAINCURSOR       <= coeff[12: 6]; 
            TXEQ_POSTCURSOR       <= coeff[17:13];
            TXEQ_NEW_COEFF[17:12] <= {1'd0, coeff[18:14]};
            TXEQ_NEW_COEFF[11: 6] <= coeff[12:7]; 
            TXEQ_NEW_COEFF[ 5: 0] <= {1'd0, coeff[5:1]}; 
            end
            
        //----------------------------------------------------------------------
        //  Hold output
        //----------------------------------------------------------------------    
        else
            begin
            TXEQ_PRECURSOR        <= TXEQ_PRECURSOR;  
            TXEQ_MAINCURSOR       <= TXEQ_MAINCURSOR; 
            TXEQ_POSTCURSOR       <= TXEQ_POSTCURSOR; 
            TXEQ_NEW_COEFF[17:12] <= TXEQ_NEW_COEFF[17:12];
            TXEQ_NEW_COEFF[11: 6] <= TXEQ_NEW_COEFF[11: 6];
            TXEQ_NEW_COEFF[ 5: 0] <= TXEQ_NEW_COEFF[ 5: 0];
            end
            
        end    
        
end



endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_gt_receiver_detect_rxterm.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//------------------------------------------------------------------------------
//  Filename     :  diablo_gt_receiver_detect_rxterm.v
//  Description  :  
//  Version      :  
//------------------------------------------------------------------------------



`timescale 1ps / 1ps



//-------------------------------------------------------------
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_gt_receiver_detect_rxterm #
(
    parameter SYNC_STAGE       = 3, 
    parameter CONSECUTIVE_CYCLE_OF_RXELECIDLE = 64
)
(
    
    //---------- Input -------------------------------------
    input               RXTERM_CLK, 
    input               RXTERM_RST_N, 
    input               RXTERM_RXELECIDLE, 
    input               RXTERM_MAC_IN_DETECT,
    
    //---------- Output ------------------------------------
    output              RXTERM_RXTERMINATION,
    output      [ 6:0]  RXTERM_FSM
);
    
    //---------- Internal Signals --------------------------
    reg                 rxelecidle_deasserted = 1'b0;
    
    //---------- Output Registers --------------------------
    reg         [ 2:0]  ctrl_fsm =  0;
    reg                 rxelecidle_int = 0;
    
    reg        [6:0]    rxelecidle_cycle_count;
    reg                 rxtermination = 0;

    wire        ctrl_fsm_not_in_solid_deassert;
    
    //---------- Control FSM ------------------------------------
    localparam          FSM_CTRL_IDLE                         = 0;
    localparam          FSM_ASSERT_AVTT                       = 1;
    localparam          FSM_CHECK_RXELECIDLE_ASSERTED         = 2; 
    localparam          FSM_CHECK_RXELECIDLE_SOLID_DEASSERT   = 3;
    localparam          FSM_ASSERT_PROG                       = 4;

    //--------------------------------------------------------------------------
    //  Synchronized Signals
    //--------------------------------------------------------------------------                                  
    wire                rxelecidle_a;
    wire                mac_in_detect_a;
    
    reg   [1:0]         rxelecidle_r;
    reg   [1:0]         mac_in_detect_r;

  xp4_usp_smsw_sync #(.WIDTH (1), .STAGE (SYNC_STAGE)) sync_rxelecidle (.CLK (RXTERM_CLK), .D (RXTERM_RXELECIDLE), .Q (rxelecidle_a));
  xp4_usp_smsw_sync #(.WIDTH (1), .STAGE (SYNC_STAGE)) sync_mac_in_detect (.CLK (RXTERM_CLK), .D (RXTERM_MAC_IN_DETECT), .Q (mac_in_detect_a));

  always @ (posedge RXTERM_CLK) 
  begin
    if (!RXTERM_RST_N) begin
      mac_in_detect_r <= 2'd3;
      rxelecidle_r <= 2'd3;
    end 
    else begin 
        rxelecidle_r <= {rxelecidle_r[0], rxelecidle_a}; 
        mac_in_detect_r <= {mac_in_detect_r[0], mac_in_detect_a};
    end
  end 
  
  always @ (posedge RXTERM_CLK) 
  begin 
    if (ctrl_fsm_not_in_solid_deassert) begin
      rxelecidle_cycle_count <= 7'd0;
    end 
    else begin
      if (!rxelecidle_a)
        rxelecidle_cycle_count <= rxelecidle_cycle_count + 7'd1;        
      else 
        rxelecidle_cycle_count <= 7'd0;
    end
  end
  
  always @(posedge RXTERM_CLK)
  begin 
    if (ctrl_fsm_not_in_solid_deassert) begin
      rxelecidle_int <= 1'b0;
    end 
    else begin
      if (rxelecidle_cycle_count > CONSECUTIVE_CYCLE_OF_RXELECIDLE)
        rxelecidle_int <= 1'b1;
      else 
        rxelecidle_int <= rxelecidle_int;
    end
  end
  
  //---------- FSM to determine when to change RX termination  --------------------
  // counter for rxelecidle. filter for consecutive #, x cycles (parameter) drive our own rxelecidle into state machine. 
  // 
  always @ (posedge RXTERM_CLK) 
  begin 
    if (!RXTERM_RST_N) begin
      ctrl_fsm   <= FSM_ASSERT_AVTT;
      rxtermination <= 1'b1;
    end
    else begin
    
      case (ctrl_fsm)
      
          //---------- Idle State ----------------------------
          FSM_CTRL_IDLE :  
            
              begin
              //----------------------------------------------
              if (!mac_in_detect_r[1]&mac_in_detect_r[0])
                  begin
                    ctrl_fsm  <= FSM_ASSERT_AVTT;
                    rxtermination <= 1'b1;
                  end
              //---------- Idle ------------------------------
              else      
                  begin
                    ctrl_fsm   <= FSM_CTRL_IDLE;
                    rxtermination <= 1'b0;
                  end
              end
              
          //---------- Assert AVTT TERMINATION ----------------
          FSM_ASSERT_AVTT :
          
              begin
                ctrl_fsm <= FSM_CHECK_RXELECIDLE_ASSERTED;
                rxtermination <= 1'b1;
              end
          
          //---------- Check RXELECIDLE is asserted --------------------
          FSM_CHECK_RXELECIDLE_ASSERTED : 
          
            begin 
              ctrl_fsm <= rxelecidle_a ? FSM_CHECK_RXELECIDLE_SOLID_DEASSERT : FSM_CHECK_RXELECIDLE_ASSERTED;
              rxtermination <= rxtermination;
            end
          
          //---------- Wait for RXELECIDELE SOLID DEASSERT and not in mac_in_detect --------------- 
          
          FSM_CHECK_RXELECIDLE_SOLID_DEASSERT:
          
              begin
                ctrl_fsm <= (rxelecidle_int&!mac_in_detect_a) ? FSM_ASSERT_PROG : FSM_CHECK_RXELECIDLE_SOLID_DEASSERT;
                rxtermination <= rxtermination;
              end

          //---------- ASSERT PROG TERMINATION -------------- 
          
          FSM_ASSERT_PROG:
          
              begin 
                ctrl_fsm <= FSM_CTRL_IDLE;
                rxtermination <= 1'b0;
              end
              
          //---------- Default State -------------------------
          default :
          
              begin      
              ctrl_fsm   <= FSM_CTRL_IDLE;
              rxtermination <= 1'b0;
              end
              
          endcase
        end
  end
  
  assign ctrl_fsm_not_in_solid_deassert = (ctrl_fsm != FSM_CHECK_RXELECIDLE_SOLID_DEASSERT);
  assign RXTERM_RXTERMINATION = rxtermination;


endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_sync_cell.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
//  Design :  PHY Wrapper
//  Module :  Synchronizer & Pipelining Cell
//--------------------------------------------------------------------------------------------------

`timescale 1ps / 1ps

//--------------------------------------------------------------------------------------------------
//  Synchronizer & Pipelining Cell 
//--------------------------------------------------------------------------------------------------
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_sync_cell #
(
    parameter integer STAGE = 3
)
(
    //-------------------------------------------------------------------------- 
    //  Input Ports
    //-------------------------------------------------------------------------- 
    input                               CLK,
    input                               D,
    
    //-------------------------------------------------------------------------- 
    //  Output Ports
    //-------------------------------------------------------------------------- 
    output                              Q
);
    //-------------------------------------------------------------------------- 
    //  Synchronized Signals
    //--------------------------------------------------------------------------  
    (* ASYNC_REG = "TRUE", SHIFT_EXTRACT = "NO" *) reg [STAGE:0] sync;                                                            



//--------------------------------------------------------------------------------------------------
//  Synchronizier
//--------------------------------------------------------------------------------------------------
always @ (posedge CLK)
begin

    sync <= {sync[(STAGE-1):0], D};
            
end   



//--------------------------------------------------------------------------------------------------
//  Generate Output
//--------------------------------------------------------------------------------------------------
assign Q = sync[STAGE];



endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_sync.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
//  Design :  PHY Wrapper
//  Module :  PHY Synchronizer & Pipelining 
//--------------------------------------------------------------------------------------------------

`timescale 1ps / 1ps

//--------------------------------------------------------------------------------------------------
//  PHY Synchronizer & Pipelining Module
//--------------------------------------------------------------------------------------------------
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_sync #
(
    parameter integer WIDTH = 1, 
    parameter integer STAGE = 3
)
(
    //-------------------------------------------------------------------------- 
    //  Input Ports
    //-------------------------------------------------------------------------- 
    input                               CLK,
    input       [WIDTH-1:0]             D,
    
    //-------------------------------------------------------------------------- 
    //  Output Ports
    //-------------------------------------------------------------------------- 
    output      [WIDTH-1:0]             Q
);                                                        



//--------------------------------------------------------------------------------------------------
//  Generate Synchronizer - Begin
//--------------------------------------------------------------------------------------------------
genvar i;

generate for (i=0; i<WIDTH; i=i+1) 

    begin : sync_vec

    //----------------------------------------------------------------------
    //  Synchronizer
    //----------------------------------------------------------------------
    xp4_usp_smsw_sync_cell #
    (
        .STAGE                          (STAGE)
    )    
    sync_cell_i
    (
        //------------------------------------------------------------------
        //  Input Ports
        //------------------------------------------------------------------
        .CLK                            (CLK),
        .D                              (D[i]),

        //------------------------------------------------------------------
        //  Output Ports
        //------------------------------------------------------------------
        .Q                              (Q[i])
    );
 
    end   
      
endgenerate 
//--------------------------------------------------------------------------------------------------
//  Generate - End
//--------------------------------------------------------------------------------------------------



endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_sys_clk_gen_ps.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//-----------------------------------------------------------------------------
//
// Project    : Ultrascale FPGA Gen4 Integrated Block for PCI Express
// File       : sys_clk_gen_ps.v
// Desc       : This file is same as sys_clk_gen.v            
// Version    : 1.0 
//-----------------------------------------------------------------------------

`timescale 1ps/1ps

module xp4_usp_smsw_sys_clk_gen_ps (sys_clk);

output	sys_clk;

reg		sys_clk;

parameter        offset = 0;
parameter        halfcycle = 500;

initial begin

	sys_clk = 0;
	#(offset);

	forever #(halfcycle) sys_clk = ~sys_clk;

end

endmodule // sys_clk_gen_ps



//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_pipe.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
/////////////////////////////////////////////////////////////////////////////

`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_pipe 
#(
     parameter           TCQ = 100
   , parameter           IMPL_TARGET = "SOFT"
   , parameter           SIM_DEVICE = "ULTRASCALE_PLUS_ES1"
   , parameter           AXISTEN_IF_EXT_512_INTFC_RAM_STYLE = "BRAM"

   , parameter           AXI4_DATA_WIDTH = 512
   , parameter           AXI4_TKEEP_WIDTH = 16
   , parameter           AXI4_CQ_TUSER_WIDTH = 183
   , parameter           AXI4_CC_TUSER_WIDTH = 81
   , parameter           AXI4_RQ_TUSER_WIDTH = 137
   , parameter           AXI4_RC_TUSER_WIDTH = 161
   , parameter           AXI4_CQ_TREADY_WIDTH = 1
   , parameter           AXI4_CC_TREADY_WIDTH = 1
   , parameter           AXI4_RQ_TREADY_WIDTH = 1
   , parameter           AXI4_RC_TREADY_WIDTH = 1

   , parameter           CRM_CORE_CLK_FREQ_500="TRUE"
   , parameter [1:0]     CRM_USER_CLK_FREQ=2'b10
   , parameter [1:0]     AXISTEN_IF_WIDTH=2'b10
   , parameter           AXISTEN_IF_EXT_512="FALSE"
   , parameter           AXISTEN_IF_EXT_512_CQ_STRADDLE="FALSE"
   , parameter           AXISTEN_IF_EXT_512_CC_STRADDLE="FALSE"
   , parameter           AXISTEN_IF_EXT_512_RQ_STRADDLE="FALSE"
   , parameter           AXISTEN_IF_EXT_512_RC_STRADDLE="FALSE"
   , parameter           AXISTEN_IF_EXT_512_RC_4TLP_STRADDLE="TRUE"
   , parameter [1:0]     AXISTEN_IF_CQ_ALIGNMENT_MODE=2'b00
   , parameter [1:0]     AXISTEN_IF_CC_ALIGNMENT_MODE=2'b00
   , parameter [1:0]     AXISTEN_IF_RQ_ALIGNMENT_MODE=2'b00
   , parameter [1:0]     AXISTEN_IF_RC_ALIGNMENT_MODE=2'b00
   , parameter           AXISTEN_IF_RC_STRADDLE="FALSE"
   , parameter           AXISTEN_IF_ENABLE_RX_MSG_INTFC="FALSE"
   , parameter [17:0]    AXISTEN_IF_ENABLE_MSG_ROUTE=18'h0
   , parameter           AXISTEN_IF_RX_PARITY_EN="TRUE"
   , parameter           AXISTEN_IF_TX_PARITY_EN="TRUE"
   , parameter           AXISTEN_IF_ENABLE_CLIENT_TAG="FALSE"
   , parameter           AXISTEN_IF_ENABLE_256_TAGS="FALSE"
   , parameter [23:0]    AXISTEN_IF_COMPL_TIMEOUT_REG0=24'hBEBC20
   , parameter [27:0]    AXISTEN_IF_COMPL_TIMEOUT_REG1=28'h2FAF080
   , parameter           AXISTEN_IF_LEGACY_MODE_ENABLE="FALSE"
   , parameter           AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK="TRUE"
   , parameter           AXISTEN_IF_MSIX_TO_RAM_PIPELINE="FALSE"
   , parameter           AXISTEN_IF_MSIX_FROM_RAM_PIPELINE="FALSE"
   , parameter           AXISTEN_IF_MSIX_RX_PARITY_EN="TRUE"
   , parameter           AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE="FALSE"
   , parameter           AXISTEN_IF_CQ_EN_POISONED_MEM_WR="FALSE"
   , parameter           AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT="FALSE"
   , parameter           AXISTEN_IF_RQ_CC_REGISTERED_TREADY="TRUE"
   , parameter [15:0]    PM_ASPML0S_TIMEOUT=16'h1500
   , parameter [31:0]    PM_L1_REENTRY_DELAY=32'h0
   , parameter [19:0]    PM_ASPML1_ENTRY_DELAY=20'h0
   , parameter           PM_ENABLE_SLOT_POWER_CAPTURE="TRUE"
   , parameter [19:0]    PM_PME_SERVICE_TIMEOUT_DELAY=20'h0
   , parameter [15:0]    PM_PME_TURNOFF_ACK_DELAY=16'h100
   , parameter           PL_UPSTREAM_FACING="TRUE"
   , parameter [4:0]     PL_LINK_CAP_MAX_LINK_WIDTH=5'b01000
   , parameter [3:0]     PL_LINK_CAP_MAX_LINK_SPEED=4'b100
   , parameter           PL_DISABLE_DC_BALANCE="FALSE"
   , parameter           PL_DISABLE_EI_INFER_IN_L0="FALSE"
   , parameter integer   PL_N_FTS=255
   , parameter           PL_DISABLE_UPCONFIG_CAPABLE="FALSE"
   , parameter           PL_DISABLE_RETRAIN_ON_FRAMING_ERROR="FALSE"
   , parameter           PL_DISABLE_RETRAIN_ON_EB_ERROR="FALSE"
   , parameter [15:0]    PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR=15'b0000000000000000
   , parameter [7:0]     PL_REPORT_ALL_PHY_ERRORS=8'b00000000
   , parameter [1:0]     PL_DISABLE_LFSR_UPDATE_ON_SKP=2'b00
   , parameter [31:0]    PL_LANE0_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE1_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE2_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE3_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE4_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE5_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE6_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE7_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE8_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE9_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE10_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE11_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE12_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE13_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE14_EQ_CONTROL=32'h3F00
   , parameter [31:0]    PL_LANE15_EQ_CONTROL=32'h3F00
   , parameter [1:0]     PL_EQ_BYPASS_PHASE23=2'b00
   , parameter [4:0]     PL_EQ_ADAPT_ITER_COUNT=5'h2
   , parameter [1:0]     PL_EQ_ADAPT_REJECT_RETRY_COUNT=2'h1
   , parameter           PL_EQ_SHORT_ADAPT_PHASE="FALSE"
   , parameter [1:0]     PL_EQ_ADAPT_DISABLE_COEFF_CHECK=2'b0
   , parameter [1:0]     PL_EQ_ADAPT_DISABLE_PRESET_CHECK=2'b0
   , parameter [7:0]     PL_EQ_DEFAULT_TX_PRESET=8'h44
   , parameter [5:0]     PL_EQ_DEFAULT_RX_PRESET_HINT=6'h33
   , parameter [1:0]     PL_EQ_RX_ADAPT_EQ_PHASE0=2'b00
   , parameter [1:0]     PL_EQ_RX_ADAPT_EQ_PHASE1=2'b00
   , parameter           PL_EQ_DISABLE_MISMATCH_CHECK="TRUE"
   , parameter [1:0]     PL_RX_L0S_EXIT_TO_RECOVERY=2'b00
   , parameter           PL_EQ_TX_8G_EQ_TS2_ENABLE="FALSE"
   , parameter           PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4="FALSE"
   , parameter           PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3="FALSE"
   , parameter           PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2="FALSE"
   , parameter           PL_DESKEW_ON_SKIP_IN_GEN12="FALSE"
   , parameter           PL_INFER_EI_DISABLE_REC_RC="FALSE"
   , parameter           PL_INFER_EI_DISABLE_REC_SPD="FALSE"
   , parameter           PL_INFER_EI_DISABLE_LPBK_ACTIVE="FALSE"
   , parameter [3:0]     PL_RX_ADAPT_TIMER_RRL_GEN3=4'h0
   , parameter [1:0]     PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS=2'b00
   , parameter [3:0]     PL_RX_ADAPT_TIMER_RRL_GEN4=4'h0
   , parameter [3:0]     PL_RX_ADAPT_TIMER_CLWS_GEN3=4'h0
   , parameter [1:0]     PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS=2'b00
   , parameter [3:0]     PL_RX_ADAPT_TIMER_CLWS_GEN4=4'h0
   , parameter           PL_DISABLE_LANE_REVERSAL="FALSE"
   , parameter           PL_CFG_STATE_ROBUSTNESS_ENABLE="TRUE"
   , parameter           PL_REDO_EQ_SOURCE_SELECT="TRUE"
   , parameter           PL_DEEMPH_SOURCE_SELECT="TRUE"
   , parameter           PL_EXIT_LOOPBACK_ON_EI_ENTRY="FALSE"
   , parameter           PL_QUIESCE_GUARANTEE_DISABLE="FALSE"
   , parameter           PL_SRIS_ENABLE="FALSE"
   , parameter [6:0]     PL_SRIS_SKPOS_GEN_SPD_VEC=7'h0
   , parameter [6:0]     PL_SRIS_SKPOS_REC_SPD_VEC=7'h0
   , parameter [1:0]     PL_SIM_FAST_LINK_TRAINING=2'h0
   , parameter [15:0]    PL_USER_SPARE=16'h0
   , parameter           LL_ACK_TIMEOUT_EN="FALSE"
   , parameter [8:0]     LL_ACK_TIMEOUT=9'h0
   , parameter integer   LL_ACK_TIMEOUT_FUNC=0
   , parameter           LL_REPLAY_TIMEOUT_EN="FALSE"
   , parameter [8:0]     LL_REPLAY_TIMEOUT=9'h0
   , parameter integer   LL_REPLAY_TIMEOUT_FUNC=0
   , parameter           LL_REPLAY_TO_RAM_PIPELINE="FALSE"
   , parameter           LL_REPLAY_FROM_RAM_PIPELINE="FALSE"
   , parameter           LL_DISABLE_SCHED_TX_NAK="FALSE"
   , parameter           LL_TX_TLP_PARITY_CHK="TRUE"
   , parameter           LL_RX_TLP_PARITY_GEN="TRUE"
   , parameter [15:0]    LL_USER_SPARE=16'h0
   , parameter           IS_SWITCH_PORT="FALSE"
   , parameter           CFG_BYPASS_MODE_ENABLE="FALSE"
   , parameter [1:0]     TL_PF_ENABLE_REG=2'h0
   , parameter [11:0]    TL_CREDITS_CD=12'h1C0
   , parameter [7:0]     TL_CREDITS_CH=8'h20
   , parameter [1:0]     TL_COMPLETION_RAM_SIZE=2'b01
   , parameter [1:0]     TL_COMPLETION_RAM_NUM_TLPS=2'b00
   , parameter [11:0]    TL_CREDITS_NPD=12'h4
   , parameter [7:0]     TL_CREDITS_NPH=8'h20
   , parameter [11:0]    TL_CREDITS_PD=12'he0
   , parameter [7:0]     TL_CREDITS_PH=8'h20
   , parameter           TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE="FALSE"
   , parameter           TL_RX_COMPLETION_TO_RAM_READ_PIPELINE="FALSE"
   , parameter           TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE="FALSE"
   , parameter           TL_POSTED_RAM_SIZE=1'b0
   , parameter           TL_RX_POSTED_TO_RAM_WRITE_PIPELINE="FALSE"
   , parameter           TL_RX_POSTED_TO_RAM_READ_PIPELINE="FALSE"
   , parameter           TL_RX_POSTED_FROM_RAM_READ_PIPELINE="FALSE"
   , parameter           TL_TX_MUX_STRICT_PRIORITY="TRUE"
   , parameter           TL_TX_TLP_STRADDLE_ENABLE="FALSE"
   , parameter           TL_TX_TLP_TERMINATE_PARITY="FALSE"
   , parameter [4:0]     TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT=5'h8
   , parameter [4:0]     TL_FC_UPDATE_MIN_INTERVAL_TIME=5'h2
   , parameter [15:0]    TL_USER_SPARE=16'h0
   , parameter [23:0]    PF0_CLASS_CODE=24'h000000
   , parameter [23:0]    PF1_CLASS_CODE=24'h000000
   , parameter [23:0]    PF2_CLASS_CODE=24'h000000
   , parameter [23:0]    PF3_CLASS_CODE=24'h000000
   , parameter [2:0]     PF0_INTERRUPT_PIN=3'h1
   , parameter [2:0]     PF1_INTERRUPT_PIN=3'h1
   , parameter [2:0]     PF2_INTERRUPT_PIN=3'h1
   , parameter [2:0]     PF3_INTERRUPT_PIN=3'h1
   , parameter [7:0]     PF0_CAPABILITY_POINTER=8'h80
   , parameter [7:0]     PF1_CAPABILITY_POINTER=8'h80
   , parameter [7:0]     PF2_CAPABILITY_POINTER=8'h80
   , parameter [7:0]     PF3_CAPABILITY_POINTER=8'h80
   , parameter [7:0]     VF0_CAPABILITY_POINTER=8'h80
   , parameter           LEGACY_CFG_EXTEND_INTERFACE_ENABLE="FALSE"
   , parameter           EXTENDED_CFG_EXTEND_INTERFACE_ENABLE="FALSE"
   , parameter           TL2CFG_IF_PARITY_CHK="TRUE"
   , parameter           HEADER_TYPE_OVERRIDE="FALSE"
   , parameter [2:0]     PF0_BAR0_CONTROL=3'b100
   , parameter [2:0]     PF1_BAR0_CONTROL=3'b100
   , parameter [2:0]     PF2_BAR0_CONTROL=3'b100
   , parameter [2:0]     PF3_BAR0_CONTROL=3'b100
   , parameter [5:0]     PF0_BAR0_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF1_BAR0_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF2_BAR0_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF3_BAR0_APERTURE_SIZE=6'b000011
   , parameter [2:0]     PF0_BAR1_CONTROL=3'b0
   , parameter [2:0]     PF1_BAR1_CONTROL=3'b0
   , parameter [2:0]     PF2_BAR1_CONTROL=3'b0
   , parameter [2:0]     PF3_BAR1_CONTROL=3'b0
   , parameter [4:0]     PF0_BAR1_APERTURE_SIZE=5'b0
   , parameter [4:0]     PF1_BAR1_APERTURE_SIZE=5'b0
   , parameter [4:0]     PF2_BAR1_APERTURE_SIZE=5'b0
   , parameter [4:0]     PF3_BAR1_APERTURE_SIZE=5'b0
   , parameter [2:0]     PF0_BAR2_CONTROL=3'b100
   , parameter [2:0]     PF1_BAR2_CONTROL=3'b100
   , parameter [2:0]     PF2_BAR2_CONTROL=3'b100
   , parameter [2:0]     PF3_BAR2_CONTROL=3'b100
   , parameter [5:0]     PF0_BAR2_APERTURE_SIZE=6'b00011
   , parameter [5:0]     PF1_BAR2_APERTURE_SIZE=6'b00011
   , parameter [5:0]     PF2_BAR2_APERTURE_SIZE=6'b00011
   , parameter [5:0]     PF3_BAR2_APERTURE_SIZE=6'b00011
   , parameter [2:0]     PF0_BAR3_CONTROL=3'b0
   , parameter [2:0]     PF1_BAR3_CONTROL=3'b0
   , parameter [2:0]     PF2_BAR3_CONTROL=3'b0
   , parameter [2:0]     PF3_BAR3_CONTROL=3'b0
   , parameter [4:0]     PF0_BAR3_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF1_BAR3_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF2_BAR3_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF3_BAR3_APERTURE_SIZE=5'b00011
   , parameter [2:0]     PF0_BAR4_CONTROL=3'b100
   , parameter [2:0]     PF1_BAR4_CONTROL=3'b100
   , parameter [2:0]     PF2_BAR4_CONTROL=3'b100
   , parameter [2:0]     PF3_BAR4_CONTROL=3'b100
   , parameter [5:0]     PF0_BAR4_APERTURE_SIZE=6'b00011
   , parameter [5:0]     PF1_BAR4_APERTURE_SIZE=6'b00011
   , parameter [5:0]     PF2_BAR4_APERTURE_SIZE=6'b00011
   , parameter [5:0]     PF3_BAR4_APERTURE_SIZE=6'b00011
   , parameter [2:0]     PF0_BAR5_CONTROL=3'b0
   , parameter [2:0]     PF1_BAR5_CONTROL=3'b0
   , parameter [2:0]     PF2_BAR5_CONTROL=3'b0
   , parameter [2:0]     PF3_BAR5_CONTROL=3'b0
   , parameter [4:0]     PF0_BAR5_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF1_BAR5_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF2_BAR5_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF3_BAR5_APERTURE_SIZE=5'b00011
   , parameter           PF0_EXPANSION_ROM_ENABLE="FALSE"
   , parameter           PF1_EXPANSION_ROM_ENABLE="FALSE"
   , parameter           PF2_EXPANSION_ROM_ENABLE="FALSE"
   , parameter           PF3_EXPANSION_ROM_ENABLE="FALSE"
   , parameter [4:0]     PF0_EXPANSION_ROM_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF1_EXPANSION_ROM_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF2_EXPANSION_ROM_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF3_EXPANSION_ROM_APERTURE_SIZE=5'b00011
   , parameter [7:0]     PF0_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF1_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF2_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF3_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     VFG0_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     VFG1_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     VFG2_PCIE_CAP_NEXTPTR=8'h0
   , parameter [7:0]     VFG3_PCIE_CAP_NEXTPTR=8'h0
   , parameter [2:0]     PF0_DEV_CAP_MAX_PAYLOAD_SIZE=3'b011
   , parameter [2:0]     PF1_DEV_CAP_MAX_PAYLOAD_SIZE=3'b011
   , parameter [2:0]     PF2_DEV_CAP_MAX_PAYLOAD_SIZE=3'b011
   , parameter [2:0]     PF3_DEV_CAP_MAX_PAYLOAD_SIZE=3'b011
   , parameter           PF0_DEV_CAP_EXT_TAG_SUPPORTED="TRUE"
   , parameter integer   PF0_DEV_CAP_ENDPOINT_L0S_LATENCY=0
   , parameter integer   PF0_DEV_CAP_ENDPOINT_L1_LATENCY=0
   , parameter           PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE="TRUE"
   , parameter integer   PF0_LINK_CAP_ASPM_SUPPORT=0
   , parameter [0:0]     PF0_LINK_CONTROL_RCB=1'b0
   , parameter           PF0_LINK_STATUS_SLOT_CLOCK_CONFIG="TRUE"
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3=7
   , parameter integer   PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3=7
   , parameter integer   PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4=7
   , parameter           PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE="TRUE"
   , parameter           PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT="TRUE"
   , parameter           PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT="TRUE"
   , parameter           PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT="TRUE"
   , parameter           PF0_DEV_CAP2_LTR_SUPPORT="TRUE"
   , parameter           PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT="FALSE"
   , parameter [1:0]     PF0_DEV_CAP2_OBFF_SUPPORT=2'b00
   , parameter           PF0_DEV_CAP2_ARI_FORWARD_ENABLE="FALSE"
   , parameter [7:0]     PF0_MSI_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF1_MSI_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF2_MSI_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF3_MSI_CAP_NEXTPTR=8'h0
   , parameter           PF0_MSI_CAP_PERVECMASKCAP="FALSE"
   , parameter           PF1_MSI_CAP_PERVECMASKCAP="FALSE"
   , parameter           PF2_MSI_CAP_PERVECMASKCAP="FALSE"
   , parameter           PF3_MSI_CAP_PERVECMASKCAP="FALSE"
   , parameter integer   PF0_MSI_CAP_MULTIMSGCAP=0
   , parameter integer   PF1_MSI_CAP_MULTIMSGCAP=0
   , parameter integer   PF2_MSI_CAP_MULTIMSGCAP=0
   , parameter integer   PF3_MSI_CAP_MULTIMSGCAP=0
   , parameter [7:0]     PF0_MSIX_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF1_MSIX_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF2_MSIX_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF3_MSIX_CAP_NEXTPTR=8'h0
   , parameter [7:0]     VFG0_MSIX_CAP_NEXTPTR=8'h0
   , parameter [7:0]     VFG1_MSIX_CAP_NEXTPTR=8'h0
   , parameter [7:0]     VFG2_MSIX_CAP_NEXTPTR=8'h0
   , parameter [7:0]     VFG3_MSIX_CAP_NEXTPTR=8'h0
   , parameter integer   PF0_MSIX_CAP_PBA_BIR=0
   , parameter integer   PF1_MSIX_CAP_PBA_BIR=0
   , parameter integer   PF2_MSIX_CAP_PBA_BIR=0
   , parameter integer   PF3_MSIX_CAP_PBA_BIR=0
   , parameter integer   VFG0_MSIX_CAP_PBA_BIR=0
   , parameter integer   VFG1_MSIX_CAP_PBA_BIR=0
   , parameter integer   VFG2_MSIX_CAP_PBA_BIR=0
   , parameter integer   VFG3_MSIX_CAP_PBA_BIR=0
   , parameter [28:0]    PF0_MSIX_CAP_PBA_OFFSET=29'h50
   , parameter [28:0]    PF1_MSIX_CAP_PBA_OFFSET=29'h50
   , parameter [28:0]    PF2_MSIX_CAP_PBA_OFFSET=29'h50
   , parameter [28:0]    PF3_MSIX_CAP_PBA_OFFSET=29'h50
   , parameter [28:0]    VFG0_MSIX_CAP_PBA_OFFSET=29'h50
   , parameter [28:0]    VFG1_MSIX_CAP_PBA_OFFSET=29'h50
   , parameter [28:0]    VFG2_MSIX_CAP_PBA_OFFSET=29'h50
   , parameter [28:0]    VFG3_MSIX_CAP_PBA_OFFSET=29'h50
   , parameter integer   PF0_MSIX_CAP_TABLE_BIR=0
   , parameter integer   PF1_MSIX_CAP_TABLE_BIR=0
   , parameter integer   PF2_MSIX_CAP_TABLE_BIR=0
   , parameter integer   PF3_MSIX_CAP_TABLE_BIR=0
   , parameter integer   VFG0_MSIX_CAP_TABLE_BIR=0
   , parameter integer   VFG1_MSIX_CAP_TABLE_BIR=0
   , parameter integer   VFG2_MSIX_CAP_TABLE_BIR=0
   , parameter integer   VFG3_MSIX_CAP_TABLE_BIR=0
   , parameter [28:0]    PF0_MSIX_CAP_TABLE_OFFSET=29'h40
   , parameter [28:0]    PF1_MSIX_CAP_TABLE_OFFSET=29'h40
   , parameter [28:0]    PF2_MSIX_CAP_TABLE_OFFSET=29'h40
   , parameter [28:0]    PF3_MSIX_CAP_TABLE_OFFSET=29'h40
   , parameter [28:0]    VFG0_MSIX_CAP_TABLE_OFFSET=29'h40
   , parameter [28:0]    VFG1_MSIX_CAP_TABLE_OFFSET=29'h40
   , parameter [28:0]    VFG2_MSIX_CAP_TABLE_OFFSET=29'h40
   , parameter [28:0]    VFG3_MSIX_CAP_TABLE_OFFSET=29'h40
   , parameter [10:0]    PF0_MSIX_CAP_TABLE_SIZE=11'h0
   , parameter [10:0]    PF1_MSIX_CAP_TABLE_SIZE=11'h0
   , parameter [10:0]    PF2_MSIX_CAP_TABLE_SIZE=11'h0
   , parameter [10:0]    PF3_MSIX_CAP_TABLE_SIZE=11'h0
   , parameter [10:0]    VFG0_MSIX_CAP_TABLE_SIZE=11'h0
   , parameter [10:0]    VFG1_MSIX_CAP_TABLE_SIZE=11'h0
   , parameter [10:0]    VFG2_MSIX_CAP_TABLE_SIZE=11'h0
   , parameter [10:0]    VFG3_MSIX_CAP_TABLE_SIZE=11'h0
   , parameter [5:0]     PF0_MSIX_VECTOR_COUNT=6'h4
   , parameter [7:0]     PF0_PM_CAP_ID=8'h1
   , parameter [7:0]     PF0_PM_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF1_PM_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF2_PM_CAP_NEXTPTR=8'h0
   , parameter [7:0]     PF3_PM_CAP_NEXTPTR=8'h0
   , parameter           PF0_PM_CAP_PMESUPPORT_D3HOT="TRUE"
   , parameter           PF0_PM_CAP_PMESUPPORT_D1="TRUE"
   , parameter           PF0_PM_CAP_PMESUPPORT_D0="TRUE"
   , parameter           PF0_PM_CAP_SUPP_D1_STATE="TRUE"
   , parameter [2:0]     PF0_PM_CAP_VER_ID=3'h3
   , parameter           PF0_PM_CSR_NOSOFTRESET="TRUE"
   , parameter           PM_ENABLE_L23_ENTRY="FALSE"
   , parameter [7:0]     DNSTREAM_LINK_NUM=8'h0
   , parameter           AUTO_FLR_RESPONSE="FALSE"
   , parameter [11:0]    PF0_DSN_CAP_NEXTPTR=12'h10C
   , parameter [11:0]    PF1_DSN_CAP_NEXTPTR=12'h10C
   , parameter [11:0]    PF2_DSN_CAP_NEXTPTR=12'h10C
   , parameter [11:0]    PF3_DSN_CAP_NEXTPTR=12'h10C
   , parameter           DSN_CAP_ENABLE="FALSE"
   , parameter [3:0]     PF0_VC_CAP_VER=4'h1
   , parameter [11:0]    PF0_VC_CAP_NEXTPTR=12'h0
   , parameter           PF0_VC_CAP_ENABLE="FALSE"
   , parameter [11:0]    PF0_SECONDARY_PCIE_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF0_AER_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF1_AER_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF2_AER_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF3_AER_CAP_NEXTPTR=12'h0
   , parameter           PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE="FALSE"
   , parameter           ARI_CAP_ENABLE="FALSE"
   , parameter [11:0]    PF0_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF1_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF2_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF3_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG0_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG1_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG2_ARI_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG3_ARI_CAP_NEXTPTR=12'h0
   , parameter [3:0]     PF0_ARI_CAP_VER=4'h1
   , parameter [7:0]     PF0_ARI_CAP_NEXT_FUNC=8'h0
   , parameter [7:0]     PF1_ARI_CAP_NEXT_FUNC=8'h0
   , parameter [7:0]     PF2_ARI_CAP_NEXT_FUNC=8'h0
   , parameter [7:0]     PF3_ARI_CAP_NEXT_FUNC=8'h0
   , parameter [11:0]    PF0_LTR_CAP_NEXTPTR=12'h0
   , parameter [3:0]     PF0_LTR_CAP_VER=4'h1
   , parameter [9:0]     PF0_LTR_CAP_MAX_SNOOP_LAT=10'h0
   , parameter [9:0]     PF0_LTR_CAP_MAX_NOSNOOP_LAT=10'h0
   , parameter           LTR_TX_MESSAGE_ON_LTR_ENABLE="FALSE"
   , parameter           LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE="FALSE"
   , parameter [9:0]     LTR_TX_MESSAGE_MINIMUM_INTERVAL=10'h250
   , parameter [3:0]     SRIOV_CAP_ENABLE=4'h0
   , parameter [11:0]    PF0_SRIOV_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF1_SRIOV_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF2_SRIOV_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF3_SRIOV_CAP_NEXTPTR=12'h0
   , parameter [3:0]     PF0_SRIOV_CAP_VER=4'h1
   , parameter [3:0]     PF1_SRIOV_CAP_VER=4'h1
   , parameter [3:0]     PF2_SRIOV_CAP_VER=4'h1
   , parameter [3:0]     PF3_SRIOV_CAP_VER=4'h1
   , parameter           PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED="FALSE"
   , parameter           PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED="FALSE"
   , parameter           PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED="FALSE"
   , parameter           PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED="FALSE"
   , parameter [15:0]    PF0_SRIOV_CAP_INITIAL_VF=16'h0
   , parameter [15:0]    PF1_SRIOV_CAP_INITIAL_VF=16'h0
   , parameter [15:0]    PF2_SRIOV_CAP_INITIAL_VF=16'h0
   , parameter [15:0]    PF3_SRIOV_CAP_INITIAL_VF=16'h0
   , parameter [15:0]    PF0_SRIOV_CAP_TOTAL_VF=16'h0
   , parameter [15:0]    PF1_SRIOV_CAP_TOTAL_VF=16'h0
   , parameter [15:0]    PF2_SRIOV_CAP_TOTAL_VF=16'h0
   , parameter [15:0]    PF3_SRIOV_CAP_TOTAL_VF=16'h0
   , parameter [15:0]    PF0_SRIOV_FUNC_DEP_LINK=16'h0
   , parameter [15:0]    PF1_SRIOV_FUNC_DEP_LINK=16'h0
   , parameter [15:0]    PF2_SRIOV_FUNC_DEP_LINK=16'h0
   , parameter [15:0]    PF3_SRIOV_FUNC_DEP_LINK=16'h0
   , parameter [15:0]    PF0_SRIOV_FIRST_VF_OFFSET=16'h0
   , parameter [15:0]    PF1_SRIOV_FIRST_VF_OFFSET=16'h0
   , parameter [15:0]    PF2_SRIOV_FIRST_VF_OFFSET=16'h0
   , parameter [15:0]    PF3_SRIOV_FIRST_VF_OFFSET=16'h0
   , parameter [15:0]    PF0_SRIOV_VF_DEVICE_ID=16'h0
   , parameter [15:0]    PF1_SRIOV_VF_DEVICE_ID=16'h0
   , parameter [15:0]    PF2_SRIOV_VF_DEVICE_ID=16'h0
   , parameter [15:0]    PF3_SRIOV_VF_DEVICE_ID=16'h0
   , parameter [31:0]    PF0_SRIOV_SUPPORTED_PAGE_SIZE=32'h0
   , parameter [31:0]    PF1_SRIOV_SUPPORTED_PAGE_SIZE=32'h0
   , parameter [31:0]    PF2_SRIOV_SUPPORTED_PAGE_SIZE=32'h0
   , parameter [31:0]    PF3_SRIOV_SUPPORTED_PAGE_SIZE=32'h0
   , parameter [2:0]     PF0_SRIOV_BAR0_CONTROL=3'b100
   , parameter [2:0]     PF1_SRIOV_BAR0_CONTROL=3'b100
   , parameter [2:0]     PF2_SRIOV_BAR0_CONTROL=3'b100
   , parameter [2:0]     PF3_SRIOV_BAR0_CONTROL=3'b100
   , parameter [5:0]     PF0_SRIOV_BAR0_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF1_SRIOV_BAR0_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF2_SRIOV_BAR0_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF3_SRIOV_BAR0_APERTURE_SIZE=6'b000011
   , parameter [2:0]     PF0_SRIOV_BAR1_CONTROL=3'b0
   , parameter [2:0]     PF1_SRIOV_BAR1_CONTROL=3'b0
   , parameter [2:0]     PF2_SRIOV_BAR1_CONTROL=3'b0
   , parameter [2:0]     PF3_SRIOV_BAR1_CONTROL=3'b0
   , parameter [4:0]     PF0_SRIOV_BAR1_APERTURE_SIZE=5'b0
   , parameter [4:0]     PF1_SRIOV_BAR1_APERTURE_SIZE=5'b0
   , parameter [4:0]     PF2_SRIOV_BAR1_APERTURE_SIZE=5'b0
   , parameter [4:0]     PF3_SRIOV_BAR1_APERTURE_SIZE=5'b0
   , parameter [2:0]     PF0_SRIOV_BAR2_CONTROL=3'b100
   , parameter [2:0]     PF1_SRIOV_BAR2_CONTROL=3'b100
   , parameter [2:0]     PF2_SRIOV_BAR2_CONTROL=3'b100
   , parameter [2:0]     PF3_SRIOV_BAR2_CONTROL=3'b100
   , parameter [5:0]     PF0_SRIOV_BAR2_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF1_SRIOV_BAR2_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF2_SRIOV_BAR2_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF3_SRIOV_BAR2_APERTURE_SIZE=6'b000011
   , parameter [2:0]     PF0_SRIOV_BAR3_CONTROL=3'b0
   , parameter [2:0]     PF1_SRIOV_BAR3_CONTROL=3'b0
   , parameter [2:0]     PF2_SRIOV_BAR3_CONTROL=3'b0
   , parameter [2:0]     PF3_SRIOV_BAR3_CONTROL=3'b0
   , parameter [4:0]     PF0_SRIOV_BAR3_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF1_SRIOV_BAR3_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF2_SRIOV_BAR3_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF3_SRIOV_BAR3_APERTURE_SIZE=5'b00011
   , parameter [2:0]     PF0_SRIOV_BAR4_CONTROL=3'b100
   , parameter [2:0]     PF1_SRIOV_BAR4_CONTROL=3'b100
   , parameter [2:0]     PF2_SRIOV_BAR4_CONTROL=3'b100
   , parameter [2:0]     PF3_SRIOV_BAR4_CONTROL=3'b100
   , parameter [5:0]     PF0_SRIOV_BAR4_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF1_SRIOV_BAR4_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF2_SRIOV_BAR4_APERTURE_SIZE=6'b000011
   , parameter [5:0]     PF3_SRIOV_BAR4_APERTURE_SIZE=6'b000011
   , parameter [2:0]     PF0_SRIOV_BAR5_CONTROL=3'b0
   , parameter [2:0]     PF1_SRIOV_BAR5_CONTROL=3'b0
   , parameter [2:0]     PF2_SRIOV_BAR5_CONTROL=3'b0
   , parameter [2:0]     PF3_SRIOV_BAR5_CONTROL=3'b0
   , parameter [4:0]     PF0_SRIOV_BAR5_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF1_SRIOV_BAR5_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF2_SRIOV_BAR5_APERTURE_SIZE=5'b00011
   , parameter [4:0]     PF3_SRIOV_BAR5_APERTURE_SIZE=5'b00011
   , parameter [11:0]    PF0_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF1_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF2_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    PF3_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG0_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG1_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG2_TPHR_CAP_NEXTPTR=12'h0
   , parameter [11:0]    VFG3_TPHR_CAP_NEXTPTR=12'h0
   , parameter [3:0]     PF0_TPHR_CAP_VER=4'h1
   , parameter           PF0_TPHR_CAP_INT_VEC_MODE="TRUE"
   , parameter           PF0_TPHR_CAP_DEV_SPECIFIC_MODE="TRUE"
   , parameter [1:0]     PF0_TPHR_CAP_ST_TABLE_LOC=2'h0
   , parameter [10:0]    PF0_TPHR_CAP_ST_TABLE_SIZE=11'h0
   , parameter [2:0]     PF0_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     PF1_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     PF2_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     PF3_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     VFG0_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     VFG1_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     VFG2_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter [2:0]     VFG3_TPHR_CAP_ST_MODE_SEL=3'h0
   , parameter           PF0_TPHR_CAP_ENABLE="FALSE"
   , parameter           TPH_TO_RAM_PIPELINE="FALSE"
   , parameter           TPH_FROM_RAM_PIPELINE="FALSE"
   , parameter           MCAP_ENABLE="FALSE"
   , parameter           MCAP_CONFIGURE_OVERRIDE="FALSE"
   , parameter [11:0]    MCAP_CAP_NEXTPTR=12'h0
   , parameter [15:0]    MCAP_VSEC_ID=16'h0
   , parameter [3:0]     MCAP_VSEC_REV=4'h0
   , parameter [11:0]    MCAP_VSEC_LEN=12'h2C
   , parameter [31:0]    MCAP_FPGA_BITSTREAM_VERSION=32'h0
   , parameter           MCAP_INTERRUPT_ON_MCAP_EOS="FALSE"
   , parameter           MCAP_INTERRUPT_ON_MCAP_ERROR="FALSE"
   , parameter           MCAP_INPUT_GATE_DESIGN_SWITCH="FALSE"
   , parameter           MCAP_EOS_DESIGN_SWITCH="FALSE"
   , parameter           MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH="FALSE"
   , parameter           MCAP_GATE_IO_ENABLE_DESIGN_SWITCH="FALSE"
   , parameter [31:0]    SIM_JTAG_IDCODE=32'h0
   , parameter [7:0]     DEBUG_AXIST_DISABLE_FEATURE_BIT=8'h0
   , parameter           DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS="FALSE"
   , parameter           DEBUG_TL_DISABLE_FC_TIMEOUT="FALSE"
   , parameter           DEBUG_PL_DISABLE_SCRAMBLING="FALSE"
   , parameter           DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL ="FALSE"
   , parameter           DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW ="FALSE"
   , parameter           DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR="FALSE"
   , parameter           DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR="FALSE"
   , parameter           DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR="FALSE"
   , parameter           DEBUG_PL_SIM_RESET_LFSR="FALSE"
   , parameter [15:0]    DEBUG_PL_SPARE=16'h0
   , parameter [15:0]    DEBUG_LL_SPARE=16'h0
   , parameter [15:0]    DEBUG_TL_SPARE=16'h0
   , parameter [15:0]    DEBUG_AXI4ST_SPARE=16'h0
   , parameter [15:0]    DEBUG_CFG_SPARE=16'h0
   , parameter [3:0]     DEBUG_CAR_SPARE=4'h0
   , parameter           TEST_MODE_PIN_CHAR="FALSE"
   , parameter           SPARE_BIT0="FALSE"
   , parameter           SPARE_BIT1=1'b0
   , parameter           SPARE_BIT2=1'b0
   , parameter           SPARE_BIT3="FALSE"
   , parameter           SPARE_BIT4=1'b0
   , parameter           SPARE_BIT5=1'b0
   , parameter           SPARE_BIT6=1'b0
   , parameter           SPARE_BIT7=1'b0
   , parameter           SPARE_BIT8=1'b0
   , parameter [7:0]     SPARE_BYTE0=8'h0
   , parameter [7:0]     SPARE_BYTE1=8'h0
   , parameter [7:0]     SPARE_BYTE2=8'h0
   , parameter [7:0]     SPARE_BYTE3=8'h0
   , parameter [31:0]    SPARE_WORD0=32'h0
   , parameter [31:0]    SPARE_WORD1=32'h0
   , parameter [31:0]    SPARE_WORD2=32'h0
   , parameter [31:0]    SPARE_WORD3=32'h0
  ) (
    input  wire [1:0]     pipe_rx00_char_is_k
   ,input  wire [1:0]     pipe_rx01_char_is_k
   ,input  wire [1:0]     pipe_rx02_char_is_k
   ,input  wire [1:0]     pipe_rx03_char_is_k
   ,input  wire [1:0]     pipe_rx04_char_is_k
   ,input  wire [1:0]     pipe_rx05_char_is_k
   ,input  wire [1:0]     pipe_rx06_char_is_k
   ,input  wire [1:0]     pipe_rx07_char_is_k
   ,input  wire [1:0]     pipe_rx08_char_is_k
   ,input  wire [1:0]     pipe_rx09_char_is_k
   ,input  wire [1:0]     pipe_rx10_char_is_k
   ,input  wire [1:0]     pipe_rx11_char_is_k
   ,input  wire [1:0]     pipe_rx12_char_is_k
   ,input  wire [1:0]     pipe_rx13_char_is_k
   ,input  wire [1:0]     pipe_rx14_char_is_k
   ,input  wire [1:0]     pipe_rx15_char_is_k
   ,input  wire           pipe_rx00_valid
   ,input  wire           pipe_rx01_valid
   ,input  wire           pipe_rx02_valid
   ,input  wire           pipe_rx03_valid
   ,input  wire           pipe_rx04_valid
   ,input  wire           pipe_rx05_valid
   ,input  wire           pipe_rx06_valid
   ,input  wire           pipe_rx07_valid
   ,input  wire           pipe_rx08_valid
   ,input  wire           pipe_rx09_valid
   ,input  wire           pipe_rx10_valid
   ,input  wire           pipe_rx11_valid
   ,input  wire           pipe_rx12_valid
   ,input  wire           pipe_rx13_valid
   ,input  wire           pipe_rx14_valid
   ,input  wire           pipe_rx15_valid
   ,input  wire [31:0]    pipe_rx00_data
   ,input  wire [31:0]    pipe_rx01_data
   ,input  wire [31:0]    pipe_rx02_data
   ,input  wire [31:0]    pipe_rx03_data
   ,input  wire [31:0]    pipe_rx04_data
   ,input  wire [31:0]    pipe_rx05_data
   ,input  wire [31:0]    pipe_rx06_data
   ,input  wire [31:0]    pipe_rx07_data
   ,input  wire [31:0]    pipe_rx08_data
   ,input  wire [31:0]    pipe_rx09_data
   ,input  wire [31:0]    pipe_rx10_data
   ,input  wire [31:0]    pipe_rx11_data
   ,input  wire [31:0]    pipe_rx12_data
   ,input  wire [31:0]    pipe_rx13_data
   ,input  wire [31:0]    pipe_rx14_data
   ,input  wire [31:0]    pipe_rx15_data
   ,output wire           pipe_rx00_polarity
   ,output wire           pipe_rx01_polarity
   ,output wire           pipe_rx02_polarity
   ,output wire           pipe_rx03_polarity
   ,output wire           pipe_rx04_polarity
   ,output wire           pipe_rx05_polarity
   ,output wire           pipe_rx06_polarity
   ,output wire           pipe_rx07_polarity
   ,output wire           pipe_rx08_polarity
   ,output wire           pipe_rx09_polarity
   ,output wire           pipe_rx10_polarity
   ,output wire           pipe_rx11_polarity
   ,output wire           pipe_rx12_polarity
   ,output wire           pipe_rx13_polarity
   ,output wire           pipe_rx14_polarity
   ,output wire           pipe_rx15_polarity
   ,input  wire [2:0]     pipe_rx00_status
   ,input  wire [2:0]     pipe_rx01_status
   ,input  wire [2:0]     pipe_rx02_status
   ,input  wire [2:0]     pipe_rx03_status
   ,input  wire [2:0]     pipe_rx04_status
   ,input  wire [2:0]     pipe_rx05_status
   ,input  wire [2:0]     pipe_rx06_status
   ,input  wire [2:0]     pipe_rx07_status
   ,input  wire [2:0]     pipe_rx08_status
   ,input  wire [2:0]     pipe_rx09_status
   ,input  wire [2:0]     pipe_rx10_status
   ,input  wire [2:0]     pipe_rx11_status
   ,input  wire [2:0]     pipe_rx12_status
   ,input  wire [2:0]     pipe_rx13_status
   ,input  wire [2:0]     pipe_rx14_status
   ,input  wire [2:0]     pipe_rx15_status
   ,input  wire           pipe_rx00_phy_status
   ,input  wire           pipe_rx01_phy_status
   ,input  wire           pipe_rx02_phy_status
   ,input  wire           pipe_rx03_phy_status
   ,input  wire           pipe_rx04_phy_status
   ,input  wire           pipe_rx05_phy_status
   ,input  wire           pipe_rx06_phy_status
   ,input  wire           pipe_rx07_phy_status
   ,input  wire           pipe_rx08_phy_status
   ,input  wire           pipe_rx09_phy_status
   ,input  wire           pipe_rx10_phy_status
   ,input  wire           pipe_rx11_phy_status
   ,input  wire           pipe_rx12_phy_status
   ,input  wire           pipe_rx13_phy_status
   ,input  wire           pipe_rx14_phy_status
   ,input  wire           pipe_rx15_phy_status
   ,input  wire           pipe_rx00_elec_idle
   ,input  wire           pipe_rx01_elec_idle
   ,input  wire           pipe_rx02_elec_idle
   ,input  wire           pipe_rx03_elec_idle
   ,input  wire           pipe_rx04_elec_idle
   ,input  wire           pipe_rx05_elec_idle
   ,input  wire           pipe_rx06_elec_idle
   ,input  wire           pipe_rx07_elec_idle
   ,input  wire           pipe_rx08_elec_idle
   ,input  wire           pipe_rx09_elec_idle
   ,input  wire           pipe_rx10_elec_idle
   ,input  wire           pipe_rx11_elec_idle
   ,input  wire           pipe_rx12_elec_idle
   ,input  wire           pipe_rx13_elec_idle
   ,input  wire           pipe_rx14_elec_idle
   ,input  wire           pipe_rx15_elec_idle
   ,input  wire           pipe_rx00_data_valid
   ,input  wire           pipe_rx01_data_valid
   ,input  wire           pipe_rx02_data_valid
   ,input  wire           pipe_rx03_data_valid
   ,input  wire           pipe_rx04_data_valid
   ,input  wire           pipe_rx05_data_valid
   ,input  wire           pipe_rx06_data_valid
   ,input  wire           pipe_rx07_data_valid
   ,input  wire           pipe_rx08_data_valid
   ,input  wire           pipe_rx09_data_valid
   ,input  wire           pipe_rx10_data_valid
   ,input  wire           pipe_rx11_data_valid
   ,input  wire           pipe_rx12_data_valid
   ,input  wire           pipe_rx13_data_valid
   ,input  wire           pipe_rx14_data_valid
   ,input  wire           pipe_rx15_data_valid
   ,input  wire [1:0]     pipe_rx00_start_block
   ,input  wire [1:0]     pipe_rx01_start_block
   ,input  wire [1:0]     pipe_rx02_start_block
   ,input  wire [1:0]     pipe_rx03_start_block
   ,input  wire [1:0]     pipe_rx04_start_block
   ,input  wire [1:0]     pipe_rx05_start_block
   ,input  wire [1:0]     pipe_rx06_start_block
   ,input  wire [1:0]     pipe_rx07_start_block
   ,input  wire [1:0]     pipe_rx08_start_block
   ,input  wire [1:0]     pipe_rx09_start_block
   ,input  wire [1:0]     pipe_rx10_start_block
   ,input  wire [1:0]     pipe_rx11_start_block
   ,input  wire [1:0]     pipe_rx12_start_block
   ,input  wire [1:0]     pipe_rx13_start_block
   ,input  wire [1:0]     pipe_rx14_start_block
   ,input  wire [1:0]     pipe_rx15_start_block
   ,input  wire [1:0]     pipe_rx00_sync_header
   ,input  wire [1:0]     pipe_rx01_sync_header
   ,input  wire [1:0]     pipe_rx02_sync_header
   ,input  wire [1:0]     pipe_rx03_sync_header
   ,input  wire [1:0]     pipe_rx04_sync_header
   ,input  wire [1:0]     pipe_rx05_sync_header
   ,input  wire [1:0]     pipe_rx06_sync_header
   ,input  wire [1:0]     pipe_rx07_sync_header
   ,input  wire [1:0]     pipe_rx08_sync_header
   ,input  wire [1:0]     pipe_rx09_sync_header
   ,input  wire [1:0]     pipe_rx10_sync_header
   ,input  wire [1:0]     pipe_rx11_sync_header
   ,input  wire [1:0]     pipe_rx12_sync_header
   ,input  wire [1:0]     pipe_rx13_sync_header
   ,input  wire [1:0]     pipe_rx14_sync_header
   ,input  wire [1:0]     pipe_rx15_sync_header
   ,output wire           pipe_tx00_compliance
   ,output wire           pipe_tx01_compliance
   ,output wire           pipe_tx02_compliance
   ,output wire           pipe_tx03_compliance
   ,output wire           pipe_tx04_compliance
   ,output wire           pipe_tx05_compliance
   ,output wire           pipe_tx06_compliance
   ,output wire           pipe_tx07_compliance
   ,output wire           pipe_tx08_compliance
   ,output wire           pipe_tx09_compliance
   ,output wire           pipe_tx10_compliance
   ,output wire           pipe_tx11_compliance
   ,output wire           pipe_tx12_compliance
   ,output wire           pipe_tx13_compliance
   ,output wire           pipe_tx14_compliance
   ,output wire           pipe_tx15_compliance
   ,output wire [1:0]     pipe_tx00_char_is_k
   ,output wire [1:0]     pipe_tx01_char_is_k
   ,output wire [1:0]     pipe_tx02_char_is_k
   ,output wire [1:0]     pipe_tx03_char_is_k
   ,output wire [1:0]     pipe_tx04_char_is_k
   ,output wire [1:0]     pipe_tx05_char_is_k
   ,output wire [1:0]     pipe_tx06_char_is_k
   ,output wire [1:0]     pipe_tx07_char_is_k
   ,output wire [1:0]     pipe_tx08_char_is_k
   ,output wire [1:0]     pipe_tx09_char_is_k
   ,output wire [1:0]     pipe_tx10_char_is_k
   ,output wire [1:0]     pipe_tx11_char_is_k
   ,output wire [1:0]     pipe_tx12_char_is_k
   ,output wire [1:0]     pipe_tx13_char_is_k
   ,output wire [1:0]     pipe_tx14_char_is_k
   ,output wire [1:0]     pipe_tx15_char_is_k
   ,output wire [31:0]    pipe_tx00_data
   ,output wire [31:0]    pipe_tx01_data
   ,output wire [31:0]    pipe_tx02_data
   ,output wire [31:0]    pipe_tx03_data
   ,output wire [31:0]    pipe_tx04_data
   ,output wire [31:0]    pipe_tx05_data
   ,output wire [31:0]    pipe_tx06_data
   ,output wire [31:0]    pipe_tx07_data
   ,output wire [31:0]    pipe_tx08_data
   ,output wire [31:0]    pipe_tx09_data
   ,output wire [31:0]    pipe_tx10_data
   ,output wire [31:0]    pipe_tx11_data
   ,output wire [31:0]    pipe_tx12_data
   ,output wire [31:0]    pipe_tx13_data
   ,output wire [31:0]    pipe_tx14_data
   ,output wire [31:0]    pipe_tx15_data
   ,output wire           pipe_tx00_elec_idle
   ,output wire           pipe_tx01_elec_idle
   ,output wire           pipe_tx02_elec_idle
   ,output wire           pipe_tx03_elec_idle
   ,output wire           pipe_tx04_elec_idle
   ,output wire           pipe_tx05_elec_idle
   ,output wire           pipe_tx06_elec_idle
   ,output wire           pipe_tx07_elec_idle
   ,output wire           pipe_tx08_elec_idle
   ,output wire           pipe_tx09_elec_idle
   ,output wire           pipe_tx10_elec_idle
   ,output wire           pipe_tx11_elec_idle
   ,output wire           pipe_tx12_elec_idle
   ,output wire           pipe_tx13_elec_idle
   ,output wire           pipe_tx14_elec_idle
   ,output wire           pipe_tx15_elec_idle
   ,output wire [1:0]     pipe_tx00_powerdown
   ,output wire [1:0]     pipe_tx01_powerdown
   ,output wire [1:0]     pipe_tx02_powerdown
   ,output wire [1:0]     pipe_tx03_powerdown
   ,output wire [1:0]     pipe_tx04_powerdown
   ,output wire [1:0]     pipe_tx05_powerdown
   ,output wire [1:0]     pipe_tx06_powerdown
   ,output wire [1:0]     pipe_tx07_powerdown
   ,output wire [1:0]     pipe_tx08_powerdown
   ,output wire [1:0]     pipe_tx09_powerdown
   ,output wire [1:0]     pipe_tx10_powerdown
   ,output wire [1:0]     pipe_tx11_powerdown
   ,output wire [1:0]     pipe_tx12_powerdown
   ,output wire [1:0]     pipe_tx13_powerdown
   ,output wire [1:0]     pipe_tx14_powerdown
   ,output wire [1:0]     pipe_tx15_powerdown
   ,output wire           pipe_tx00_data_valid
   ,output wire           pipe_tx01_data_valid
   ,output wire           pipe_tx02_data_valid
   ,output wire           pipe_tx03_data_valid
   ,output wire           pipe_tx04_data_valid
   ,output wire           pipe_tx05_data_valid
   ,output wire           pipe_tx06_data_valid
   ,output wire           pipe_tx07_data_valid
   ,output wire           pipe_tx08_data_valid
   ,output wire           pipe_tx09_data_valid
   ,output wire           pipe_tx10_data_valid
   ,output wire           pipe_tx11_data_valid
   ,output wire           pipe_tx12_data_valid
   ,output wire           pipe_tx13_data_valid
   ,output wire           pipe_tx14_data_valid
   ,output wire           pipe_tx15_data_valid
   ,output wire           pipe_tx00_start_block
   ,output wire           pipe_tx01_start_block
   ,output wire           pipe_tx02_start_block
   ,output wire           pipe_tx03_start_block
   ,output wire           pipe_tx04_start_block
   ,output wire           pipe_tx05_start_block
   ,output wire           pipe_tx06_start_block
   ,output wire           pipe_tx07_start_block
   ,output wire           pipe_tx08_start_block
   ,output wire           pipe_tx09_start_block
   ,output wire           pipe_tx10_start_block
   ,output wire           pipe_tx11_start_block
   ,output wire           pipe_tx12_start_block
   ,output wire           pipe_tx13_start_block
   ,output wire           pipe_tx14_start_block
   ,output wire           pipe_tx15_start_block
   ,output wire [1:0]     pipe_tx00_sync_header
   ,output wire [1:0]     pipe_tx01_sync_header
   ,output wire [1:0]     pipe_tx02_sync_header
   ,output wire [1:0]     pipe_tx03_sync_header
   ,output wire [1:0]     pipe_tx04_sync_header
   ,output wire [1:0]     pipe_tx05_sync_header
   ,output wire [1:0]     pipe_tx06_sync_header
   ,output wire [1:0]     pipe_tx07_sync_header
   ,output wire [1:0]     pipe_tx08_sync_header
   ,output wire [1:0]     pipe_tx09_sync_header
   ,output wire [1:0]     pipe_tx10_sync_header
   ,output wire [1:0]     pipe_tx11_sync_header
   ,output wire [1:0]     pipe_tx12_sync_header
   ,output wire [1:0]     pipe_tx13_sync_header
   ,output wire [1:0]     pipe_tx14_sync_header
   ,output wire [1:0]     pipe_tx15_sync_header
   ,output wire [1:0]     pipe_rx00_eq_control
   ,output wire [1:0]     pipe_rx01_eq_control
   ,output wire [1:0]     pipe_rx02_eq_control
   ,output wire [1:0]     pipe_rx03_eq_control
   ,output wire [1:0]     pipe_rx04_eq_control
   ,output wire [1:0]     pipe_rx05_eq_control
   ,output wire [1:0]     pipe_rx06_eq_control
   ,output wire [1:0]     pipe_rx07_eq_control
   ,output wire [1:0]     pipe_rx08_eq_control
   ,output wire [1:0]     pipe_rx09_eq_control
   ,output wire [1:0]     pipe_rx10_eq_control
   ,output wire [1:0]     pipe_rx11_eq_control
   ,output wire [1:0]     pipe_rx12_eq_control
   ,output wire [1:0]     pipe_rx13_eq_control
   ,output wire [1:0]     pipe_rx14_eq_control
   ,output wire [1:0]     pipe_rx15_eq_control
   ,input  wire           pipe_rx00_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx01_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx02_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx03_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx04_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx05_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx06_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx07_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx08_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx09_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx10_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx11_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx12_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx13_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx14_eq_lp_lf_fs_sel
   ,input  wire           pipe_rx15_eq_lp_lf_fs_sel
   ,input  wire [17:0]    pipe_rx00_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx01_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx02_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx03_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx04_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx05_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx06_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx07_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx08_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx09_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx10_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx11_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx12_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx13_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx14_eq_lp_new_tx_coeff_or_preset
   ,input  wire [17:0]    pipe_rx15_eq_lp_new_tx_coeff_or_preset
   ,input  wire           pipe_rx00_eq_lp_adapt_done
   ,input  wire           pipe_rx01_eq_lp_adapt_done
   ,input  wire           pipe_rx02_eq_lp_adapt_done
   ,input  wire           pipe_rx03_eq_lp_adapt_done
   ,input  wire           pipe_rx04_eq_lp_adapt_done
   ,input  wire           pipe_rx05_eq_lp_adapt_done
   ,input  wire           pipe_rx06_eq_lp_adapt_done
   ,input  wire           pipe_rx07_eq_lp_adapt_done
   ,input  wire           pipe_rx08_eq_lp_adapt_done
   ,input  wire           pipe_rx09_eq_lp_adapt_done
   ,input  wire           pipe_rx10_eq_lp_adapt_done
   ,input  wire           pipe_rx11_eq_lp_adapt_done
   ,input  wire           pipe_rx12_eq_lp_adapt_done
   ,input  wire           pipe_rx13_eq_lp_adapt_done
   ,input  wire           pipe_rx14_eq_lp_adapt_done
   ,input  wire           pipe_rx15_eq_lp_adapt_done
   ,input  wire           pipe_rx00_eq_done
   ,input  wire           pipe_rx01_eq_done
   ,input  wire           pipe_rx02_eq_done
   ,input  wire           pipe_rx03_eq_done
   ,input  wire           pipe_rx04_eq_done
   ,input  wire           pipe_rx05_eq_done
   ,input  wire           pipe_rx06_eq_done
   ,input  wire           pipe_rx07_eq_done
   ,input  wire           pipe_rx08_eq_done
   ,input  wire           pipe_rx09_eq_done
   ,input  wire           pipe_rx10_eq_done
   ,input  wire           pipe_rx11_eq_done
   ,input  wire           pipe_rx12_eq_done
   ,input  wire           pipe_rx13_eq_done
   ,input  wire           pipe_rx14_eq_done
   ,input  wire           pipe_rx15_eq_done
   ,output wire [1:0]     pipe_tx00_eq_control
   ,output wire [1:0]     pipe_tx01_eq_control
   ,output wire [1:0]     pipe_tx02_eq_control
   ,output wire [1:0]     pipe_tx03_eq_control
   ,output wire [1:0]     pipe_tx04_eq_control
   ,output wire [1:0]     pipe_tx05_eq_control
   ,output wire [1:0]     pipe_tx06_eq_control
   ,output wire [1:0]     pipe_tx07_eq_control
   ,output wire [1:0]     pipe_tx08_eq_control
   ,output wire [1:0]     pipe_tx09_eq_control
   ,output wire [1:0]     pipe_tx10_eq_control
   ,output wire [1:0]     pipe_tx11_eq_control
   ,output wire [1:0]     pipe_tx12_eq_control
   ,output wire [1:0]     pipe_tx13_eq_control
   ,output wire [1:0]     pipe_tx14_eq_control
   ,output wire [1:0]     pipe_tx15_eq_control
   ,output wire [5:0]     pipe_tx00_eq_deemph
   ,output wire [5:0]     pipe_tx01_eq_deemph
   ,output wire [5:0]     pipe_tx02_eq_deemph
   ,output wire [5:0]     pipe_tx03_eq_deemph
   ,output wire [5:0]     pipe_tx04_eq_deemph
   ,output wire [5:0]     pipe_tx05_eq_deemph
   ,output wire [5:0]     pipe_tx06_eq_deemph
   ,output wire [5:0]     pipe_tx07_eq_deemph
   ,output wire [5:0]     pipe_tx08_eq_deemph
   ,output wire [5:0]     pipe_tx09_eq_deemph
   ,output wire [5:0]     pipe_tx10_eq_deemph
   ,output wire [5:0]     pipe_tx11_eq_deemph
   ,output wire [5:0]     pipe_tx12_eq_deemph
   ,output wire [5:0]     pipe_tx13_eq_deemph
   ,output wire [5:0]     pipe_tx14_eq_deemph
   ,output wire [5:0]     pipe_tx15_eq_deemph
   ,input  wire [17:0]    pipe_tx00_eq_coeff
   ,input  wire [17:0]    pipe_tx01_eq_coeff
   ,input  wire [17:0]    pipe_tx02_eq_coeff
   ,input  wire [17:0]    pipe_tx03_eq_coeff
   ,input  wire [17:0]    pipe_tx04_eq_coeff
   ,input  wire [17:0]    pipe_tx05_eq_coeff
   ,input  wire [17:0]    pipe_tx06_eq_coeff
   ,input  wire [17:0]    pipe_tx07_eq_coeff
   ,input  wire [17:0]    pipe_tx08_eq_coeff
   ,input  wire [17:0]    pipe_tx09_eq_coeff
   ,input  wire [17:0]    pipe_tx10_eq_coeff
   ,input  wire [17:0]    pipe_tx11_eq_coeff
   ,input  wire [17:0]    pipe_tx12_eq_coeff
   ,input  wire [17:0]    pipe_tx13_eq_coeff
   ,input  wire [17:0]    pipe_tx14_eq_coeff
   ,input  wire [17:0]    pipe_tx15_eq_coeff
   ,input  wire           pipe_tx00_eq_done
   ,input  wire           pipe_tx01_eq_done
   ,input  wire           pipe_tx02_eq_done
   ,input  wire           pipe_tx03_eq_done
   ,input  wire           pipe_tx04_eq_done
   ,input  wire           pipe_tx05_eq_done
   ,input  wire           pipe_tx06_eq_done
   ,input  wire           pipe_tx07_eq_done
   ,input  wire           pipe_tx08_eq_done
   ,input  wire           pipe_tx09_eq_done
   ,input  wire           pipe_tx10_eq_done
   ,input  wire           pipe_tx11_eq_done
   ,input  wire           pipe_tx12_eq_done
   ,input  wire           pipe_tx13_eq_done
   ,input  wire           pipe_tx14_eq_done
   ,input  wire           pipe_tx15_eq_done
   ,output wire [3:0]     pipe_rx_eq_lp_tx_preset
   ,output wire [5:0]     pipe_rx_eq_lp_lf_fs
   ,output wire           pipe_tx_rcvr_det
   ,output wire [1:0]     pipe_tx_rate
   ,output wire           pipe_tx_deemph
   ,output wire [2:0]     pipe_tx_margin
   ,output wire           pipe_tx_swing
   ,output wire           pipe_tx_reset
   ,input  wire [5:0]     pipe_eq_fs
   ,input  wire [5:0]     pipe_eq_lf
   ,input  wire           pl_gen2_upstream_prefer_deemph
   ,output wire           pl_eq_in_progress
   ,output wire [1:0]     pl_eq_phase
   ,input  wire           pl_eq_reset_eieos_count
   ,input  wire           pl_redo_eq
   ,input  wire           pl_redo_eq_speed
   ,output wire           pl_eq_mismatch
   ,output wire           pl_redo_eq_pending
   ,output wire [AXI4_DATA_WIDTH-1:0] m_axis_cq_tdata
   ,input  wire [AXI4_DATA_WIDTH-1:0] s_axis_cc_tdata
   ,input  wire [AXI4_DATA_WIDTH-1:0] s_axis_rq_tdata
   ,output wire [AXI4_DATA_WIDTH-1:0] m_axis_rc_tdata
   ,output wire [AXI4_CQ_TUSER_WIDTH-1:0] m_axis_cq_tuser
   ,input  wire [AXI4_CC_TUSER_WIDTH-1:0] s_axis_cc_tuser
   ,output wire           m_axis_cq_tlast
   ,input  wire           s_axis_rq_tlast
   ,output wire           m_axis_rc_tlast
   ,input  wire           s_axis_cc_tlast
   ,input  wire [1:0]     pcie_cq_np_req
   ,output wire [5:0]     pcie_cq_np_req_count
   ,input  wire [AXI4_RQ_TUSER_WIDTH-1:0] s_axis_rq_tuser
   ,output wire [AXI4_RC_TUSER_WIDTH-1:0] m_axis_rc_tuser
   ,output wire [AXI4_TKEEP_WIDTH-1:0] m_axis_cq_tkeep
   ,input  wire [AXI4_TKEEP_WIDTH-1:0] s_axis_cc_tkeep
   ,input  wire [AXI4_TKEEP_WIDTH-1:0] s_axis_rq_tkeep
   ,output wire [AXI4_TKEEP_WIDTH-1:0] m_axis_rc_tkeep
   ,output wire           m_axis_cq_tvalid
   ,input  wire           s_axis_cc_tvalid
   ,input  wire           s_axis_rq_tvalid
   ,output wire           m_axis_rc_tvalid
   ,input  wire [AXI4_CQ_TREADY_WIDTH-1:0] m_axis_cq_tready
   ,output wire [AXI4_CC_TREADY_WIDTH-1:0] s_axis_cc_tready
   ,output wire [AXI4_RQ_TREADY_WIDTH-1:0] s_axis_rq_tready
   ,input  wire [AXI4_RC_TREADY_WIDTH-1:0] m_axis_rc_tready
   ,output wire [5:0]     pcie_rq_seq_num0
   ,output wire           pcie_rq_seq_num_vld0
   ,output wire [5:0]     pcie_rq_seq_num1
   ,output wire           pcie_rq_seq_num_vld1
   ,output wire [7:0]     pcie_rq_tag0
   ,output wire           pcie_rq_tag_vld0
   ,output wire [7:0]     pcie_rq_tag1
   ,output wire           pcie_rq_tag_vld1
   ,output wire [3:0]     pcie_tfc_nph_av
   ,output wire [3:0]     pcie_tfc_npd_av
   ,output wire [3:0]     pcie_rq_tag_av
   ,output wire [7:0]     axi_user_out
   ,input  wire [7:0]     axi_user_in
   ,input  wire [9:0]     cfg_mgmt_addr
   ,input  wire [7:0]     cfg_mgmt_function_number
   ,input  wire           cfg_mgmt_write
   ,input  wire [31:0]    cfg_mgmt_write_data
   ,input  wire [3:0]     cfg_mgmt_byte_enable
   ,input  wire           cfg_mgmt_read
   ,output wire [31:0]    cfg_mgmt_read_data
   ,output wire           cfg_mgmt_read_write_done
   ,input  wire           cfg_mgmt_debug_access
   ,output wire           cfg_phy_link_down
   ,output wire [1:0]     cfg_phy_link_status
   ,output wire [2:0]     cfg_negotiated_width
   ,output wire [1:0]     cfg_current_speed
   ,output wire [1:0]     cfg_max_payload
   ,output wire [2:0]     cfg_max_read_req
   ,output wire [15:0]    cfg_function_status
   ,output wire [11:0]    cfg_function_power_state
   ,output wire [1:0]     cfg_link_power_state
   ,output wire           cfg_err_cor_out
   ,output wire           cfg_err_nonfatal_out
   ,output wire           cfg_err_fatal_out
   ,output wire           cfg_local_error_valid
   ,output wire [4:0]     cfg_local_error_out
   ,output wire           cfg_ltr_enable
   ,output wire [5:0]     cfg_ltssm_state
   ,output wire [1:0]     cfg_rx_pm_state
   ,output wire [1:0]     cfg_tx_pm_state
   ,output wire [3:0]     cfg_rcb_status
   ,output wire [1:0]     cfg_obff_enable
   ,output wire           cfg_pl_status_change
   ,output wire [3:0]     cfg_tph_requester_enable
   ,output wire [11:0]    cfg_tph_st_mode
   ,output wire           cfg_msg_received
   ,output wire [7:0]     cfg_msg_received_data
   ,output wire [4:0]     cfg_msg_received_type
   ,input  wire           cfg_msg_transmit
   ,input  wire [2:0]     cfg_msg_transmit_type
   ,input  wire [31:0]    cfg_msg_transmit_data
   ,output wire           cfg_msg_transmit_done
   ,output wire [7:0]     cfg_fc_ph
   ,output wire [11:0]    cfg_fc_pd
   ,output wire [7:0]     cfg_fc_nph
   ,output wire [11:0]    cfg_fc_npd
   ,output wire [7:0]     cfg_fc_cplh
   ,output wire [11:0]    cfg_fc_cpld
   ,input  wire [2:0]     cfg_fc_sel
   ,input  wire           cfg_hot_reset_in
   ,output wire           cfg_hot_reset_out
   ,input  wire           cfg_config_space_enable
   ,input  wire [63:0]    cfg_dsn
   ,input  wire [15:0]    cfg_dev_id_pf0
   ,input  wire [15:0]    cfg_dev_id_pf1
   ,input  wire [15:0]    cfg_dev_id_pf2
   ,input  wire [15:0]    cfg_dev_id_pf3
   ,input  wire [15:0]    cfg_vend_id
   ,input  wire [7:0]     cfg_rev_id_pf0
   ,input  wire [7:0]     cfg_rev_id_pf1
   ,input  wire [7:0]     cfg_rev_id_pf2
   ,input  wire [7:0]     cfg_rev_id_pf3
   ,input  wire [15:0]    cfg_subsys_id_pf0
   ,input  wire [15:0]    cfg_subsys_id_pf1
   ,input  wire [15:0]    cfg_subsys_id_pf2
   ,input  wire [15:0]    cfg_subsys_id_pf3
   ,input  wire [15:0]    cfg_subsys_vend_id
   ,input  wire [7:0]     cfg_ds_port_number
   ,input  wire [7:0]     cfg_ds_bus_number
   ,input  wire [4:0]     cfg_ds_device_number
   ,input  wire [2:0]     cfg_ds_function_number
   ,output wire [7:0]     cfg_bus_number
   ,input  wire           cfg_power_state_change_ack
   ,output wire           cfg_power_state_change_interrupt
   ,input  wire           cfg_err_cor_in
   ,input  wire           cfg_err_uncor_in
   ,input  wire [3:0]     cfg_flr_done
   ,output wire [3:0]     cfg_flr_in_process
   ,input  wire           cfg_req_pm_transition_l23_ready
   ,input  wire           cfg_link_training_enable
   ,input  wire [3:0]     cfg_interrupt_int
   ,output wire           cfg_interrupt_sent
   ,input  wire [3:0]     cfg_interrupt_pending
   ,output wire [3:0]     cfg_interrupt_msi_enable
   ,input  wire [31:0]    cfg_interrupt_msi_int
   ,output wire           cfg_interrupt_msi_sent
   ,output wire           cfg_interrupt_msi_fail
   ,output wire [11:0]    cfg_interrupt_msi_mmenable
   ,input  wire [31:0]    cfg_interrupt_msi_pending_status
   ,input  wire [1:0]     cfg_interrupt_msi_pending_status_function_num
   ,input  wire           cfg_interrupt_msi_pending_status_data_enable
   ,output wire           cfg_interrupt_msi_mask_update
   ,input  wire [1:0]     cfg_interrupt_msi_select
   ,output wire [31:0]    cfg_interrupt_msi_data
   ,output wire [3:0]     cfg_interrupt_msix_enable
   ,output wire [3:0]     cfg_interrupt_msix_mask
   ,input  wire [63:0]    cfg_interrupt_msix_address
   ,input  wire [31:0]    cfg_interrupt_msix_data
   ,input  wire           cfg_interrupt_msix_int
   ,input  wire [1:0]     cfg_interrupt_msix_vec_pending
   ,output wire           cfg_interrupt_msix_vec_pending_status
   ,input  wire [2:0]     cfg_interrupt_msi_attr
   ,input  wire           cfg_interrupt_msi_tph_present
   ,input  wire [1:0]     cfg_interrupt_msi_tph_type
   ,input  wire [7:0]     cfg_interrupt_msi_tph_st_tag
   ,input  wire [7:0]     cfg_interrupt_msi_function_number
   ,output wire           cfg_ext_read_received
   ,output wire           cfg_ext_write_received
   ,output wire [9:0]     cfg_ext_register_number
   ,output wire [7:0]     cfg_ext_function_number
   ,output wire [31:0]    cfg_ext_write_data
   ,output wire [3:0]     cfg_ext_write_byte_enable
   ,input  wire [31:0]    cfg_ext_read_data
   ,input  wire           cfg_ext_read_data_valid
   ,output wire [251:0]   cfg_vf_flr_in_process
   ,input  wire [7:0]     cfg_vf_flr_func_num
   ,input  wire           cfg_vf_flr_done
   ,output wire [503:0]   cfg_vf_status
   ,output wire [755:0]   cfg_vf_power_state
   ,output wire [251:0]   cfg_vf_tph_requester_enable
   ,output wire [755:0]   cfg_vf_tph_st_mode
   ,output wire [251:0]   cfg_interrupt_msix_vf_enable
   ,output wire [251:0]   cfg_interrupt_msix_vf_mask
   ,input  wire           cfg_pm_aspm_l1_entry_reject
   ,input  wire           cfg_pm_aspm_tx_l0s_entry_disable
   ,input  wire [7:0]     user_tph_stt_func_num
   ,input  wire [5:0]     user_tph_stt_index
   ,input  wire           user_tph_stt_rd_en
   ,output wire [7:0]     user_tph_stt_rd_data
   ,input  wire [1:0]     conf_req_type
   ,input  wire [3:0]     conf_req_reg_num
   ,input  wire [31:0]    conf_req_data
   ,input  wire           conf_req_valid
   ,output wire           conf_req_ready
   ,output wire [31:0]    conf_resp_rdata
   ,output wire           conf_resp_valid
   ,output wire           conf_mcap_design_switch
   ,output wire           conf_mcap_eos
   ,output wire           conf_mcap_in_use_by_pcie
   ,input  wire           conf_mcap_request_by_conf
   ,input  wire           drp_clk
   ,input  wire           drp_en
   ,input  wire           drp_we
   ,input  wire [9:0]     drp_addr
   ,input  wire [15:0]    drp_di
   ,output wire           drp_rdy
   ,output wire [15:0]    drp_do

   ,input  wire           pipe_clk
   ,input  wire           core_clk
   ,input  wire           user_clk
   ,input  wire           user_clk2
   ,output wire           user_clk_en
   ,input  wire           mcap_clk
   ,input  wire           mcap_rst_b
   ,output wire           pcie_perst0_b
   ,output wire           pcie_perst1_b
   ,input  wire           phy_rdy 
  );

  // localparams
  
  localparam [10:0]      MSIX_CAP_TABLE_SIZE = PF0_MSIX_CAP_TABLE_SIZE +
                                               PF1_MSIX_CAP_TABLE_SIZE +
                                               PF2_MSIX_CAP_TABLE_SIZE +
                                               PF3_MSIX_CAP_TABLE_SIZE +
                                               VFG0_MSIX_CAP_TABLE_SIZE +
                                               VFG1_MSIX_CAP_TABLE_SIZE +
                                               VFG2_MSIX_CAP_TABLE_SIZE +
                                               VFG3_MSIX_CAP_TABLE_SIZE;
  localparam             MSIX_TABLE_RAM_ENABLE = AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE;


  // Resets
  
  wire                        reset_n;
  wire                        mgmt_reset_n;
  wire                        mgmt_sticky_reset_n;
  wire                        pipe_reset_n;
  wire                        user_clkgate_en;
  wire                        pipe_clkgate_en;
  wire                        user_clk_en_to_e4;
  wire                        user_clk_to_e4;
  wire                        user_clk2_to_e4;
  wire                        pipe_clk_to_e4;
  wire                        cfg_phy_link_down_wire;
  wire                        cfg_phy_link_down_user_clk;

  wire [31:0]                 pipe_tx00_data_out;
  wire [31:0]                 pipe_tx01_data_out;
  wire [31:0]                 pipe_tx02_data_out;
  wire [31:0]                 pipe_tx03_data_out;
  wire [31:0]                 pipe_tx04_data_out;
  wire [31:0]                 pipe_tx05_data_out;
  wire [31:0]                 pipe_tx06_data_out;
  wire [31:0]                 pipe_tx07_data_out;
  wire [31:0]                 pipe_tx08_data_out;
  wire [31:0]                 pipe_tx09_data_out;
  wire [31:0]                 pipe_tx10_data_out;
  wire [31:0]                 pipe_tx11_data_out;
  wire [31:0]                 pipe_tx12_data_out;
  wire [31:0]                 pipe_tx13_data_out;
  wire [31:0]                 pipe_tx14_data_out;
  wire [31:0]                 pipe_tx15_data_out;

  assign cfg_phy_link_down = cfg_phy_link_down_wire;

generate if (IMPL_TARGET=="SOFT" || IMPL_TARGET=="PROTO") begin

   // no clock gating case for soft or hard
   assign user_clk_en_to_e4  = user_clk_en;
   assign user_clk_to_e4     = user_clk;
   assign user_clk2_to_e4    = user_clk2;
   assign pipe_clk_to_e4     = pipe_clk;   

end else begin

   // clock gating case for soft or hard
   assign user_clk_en_to_e4  = user_clkgate_en;
   assign user_clk_to_e4     = 1'b0;
   assign user_clk2_to_e4    = 1'b0;
   assign pipe_clk_to_e4     = pipe_clk;   // pipe clock gating not yet included

end
endgenerate

    assign pipe_tx00_data = pipe_tx00_data_out; 
    assign pipe_tx01_data = pipe_tx01_data_out;
    assign pipe_tx02_data = pipe_tx02_data_out;
    assign pipe_tx03_data = pipe_tx03_data_out;
    assign pipe_tx04_data = pipe_tx04_data_out;
    assign pipe_tx05_data = pipe_tx05_data_out;
    assign pipe_tx06_data = pipe_tx06_data_out;
    assign pipe_tx07_data = pipe_tx07_data_out;
    assign pipe_tx08_data = pipe_tx08_data_out;
    assign pipe_tx09_data = pipe_tx09_data_out;
    assign pipe_tx10_data = pipe_tx10_data_out;
    assign pipe_tx11_data = pipe_tx11_data_out;
    assign pipe_tx12_data = pipe_tx12_data_out;
    assign pipe_tx13_data = pipe_tx13_data_out;
    assign pipe_tx14_data = pipe_tx14_data_out;
    assign pipe_tx15_data = pipe_tx15_data_out;
     
   
  // Memory Interfaces

  wire [8:0]                  mi_replay_ram_address0;
  wire [8:0]                  mi_replay_ram_address1;
  wire [127:0]                mi_replay_ram_write_data0;
  wire                        mi_replay_ram_write_enable0;
  wire [127:0]                mi_replay_ram_write_data1;
  wire                        mi_replay_ram_write_enable1;
  wire [127:0]                mi_replay_ram_read_data0;
  wire                        mi_replay_ram_read_enable0;
  wire [127:0]                mi_replay_ram_read_data1;
  wire                        mi_replay_ram_read_enable1;
  wire [5:0]                  mi_replay_ram_err_cor;
  wire [5:0]                  mi_replay_ram_err_uncor;
  wire [8:0]                  mi_rx_posted_request_ram_write_address0;
  wire [143:0]                mi_rx_posted_request_ram_write_data0;
  wire                        mi_rx_posted_request_ram_write_enable0;
  wire [8:0]                  mi_rx_posted_request_ram_write_address1;
  wire [143:0]                mi_rx_posted_request_ram_write_data1;
  wire                        mi_rx_posted_request_ram_write_enable1;
  wire [8:0]                  mi_rx_posted_request_ram_read_address0;
  wire [143:0]                mi_rx_posted_request_ram_read_data0;
  wire                        mi_rx_posted_request_ram_read_enable0;
  wire [8:0]                  mi_rx_posted_request_ram_read_address1;
  wire [143:0]                mi_rx_posted_request_ram_read_data1;
  wire                        mi_rx_posted_request_ram_read_enable1;
  wire [5:0]                  mi_rx_posted_request_ram_err_cor;
  wire [5:0]                  mi_rx_posted_request_ram_err_uncor;
  wire [8:0]                  mi_rx_completion_ram_write_address0;
  wire [143:0]                mi_rx_completion_ram_write_data0;
  wire [1:0]                  mi_rx_completion_ram_write_enable0;
  wire [8:0]                  mi_rx_completion_ram_write_address1;
  wire [143:0]                mi_rx_completion_ram_write_data1;
  wire [1:0]                  mi_rx_completion_ram_write_enable1;
  wire [8:0]                  mi_rx_completion_ram_read_address0;
  wire [143:0]                mi_rx_completion_ram_read_data0;
  wire [1:0]                  mi_rx_completion_ram_read_enable0;
  wire [8:0]                  mi_rx_completion_ram_read_address1;
  wire [143:0]                mi_rx_completion_ram_read_data1;
  wire [1:0]                  mi_rx_completion_ram_read_enable1;
  wire [11:0]                 mi_rx_completion_ram_err_cor;
  wire [11:0]                 mi_rx_completion_ram_err_uncor;
  wire [11:0]                 cfg_tph_ram_address;
  wire [35:0]                 cfg_tph_ram_write_data;
  wire [3:0]                  cfg_tph_ram_write_byte_enable;
  wire [35:0]                 cfg_tph_ram_read_data;
  wire                        cfg_tph_ram_read_enable;
  wire [12:0]                 cfg_msix_ram_address;
  wire [35:0]                 cfg_msix_ram_write_data;
  wire [3:0]                  cfg_msix_ram_write_byte_enable;
  wire [35:0]                 cfg_msix_ram_read_data;
  wire                        cfg_msix_ram_read_enable;
 
  // Driven by soft logic
  wire                        pcie_posted_req_delivered;
  wire                        pcie_cq_pipeline_empty;
  wire                        pcie_cq_np_user_credit_rcvd;
  wire [1:0]                  pcie_compl_delivered;
  wire [7:0]                  pcie_compl_delivered_tag0;
  wire [7:0]                  pcie_compl_delivered_tag1;

  // Wires from Hard Block AXI Stream Interface to Soft Bridge
  wire [255:0]                m_axis_cq_tdata_int;
  wire [87:0]                 m_axis_cq_tuser_int;
  wire                        m_axis_cq_tlast_int;
  wire [7:0]                  m_axis_cq_tkeep_int;
  wire                        m_axis_cq_tvalid_int;
        
  wire [255:0]                s_axis_cc_tdata_int;
  wire [32:0]                 s_axis_cc_tuser_int;
  wire                        s_axis_cc_tlast_int;
  wire [7:0]                  s_axis_cc_tkeep_int;
  wire                        s_axis_cc_tvalid_int;

  wire [255:0]                s_axis_rq_tdata_int;
  wire [61:0]                 s_axis_rq_tuser_int;
  wire                        s_axis_rq_tlast_int;
  wire [7:0]                  s_axis_rq_tkeep_int;
  wire                        s_axis_rq_tvalid_int;

  wire [255:0]                m_axis_rc_tdata_int;
  wire [74:0]                 m_axis_rc_tuser_int;
  wire                        m_axis_rc_tlast_int;
  wire [7:0]                  m_axis_rc_tkeep_int;
  wire                        m_axis_rc_tvalid_int;

  wire [255:0]                s_axis_cc_tdata_axi512;
  wire [32:0]                 s_axis_cc_tuser_axi512;
  wire                        s_axis_cc_tlast_axi512;
  wire [7:0]                  s_axis_cc_tkeep_axi512;
  wire                        s_axis_cc_tvalid_axi512;

  wire [255:0]                s_axis_rq_tdata_axi512;
  wire [61:0]                 s_axis_rq_tuser_axi512;
  wire                        s_axis_rq_tlast_axi512;
  wire [7:0]                  s_axis_rq_tkeep_axi512;
  wire                        s_axis_rq_tvalid_axi512;

  wire [21:0]                 m_axis_cq_tready_int;
  wire [21:0]                 m_axis_rc_tready_int;
  wire [21:0]                 m_axis_cq_tready_axi512;
  wire [21:0]                 m_axis_rc_tready_axi512;
  wire [3:0]                  s_axis_cc_tready_int;
  wire                        s_axis_cc_tready_axi512;
  wire [3:0]                  s_axis_rq_tready_int;
  wire                        s_axis_rq_tready_axi512;

  wire [5:0]                  pcie_cq_np_req_count_int;
  wire [5:0]                  pcie_cq_np_req_count_axi512;

  wire                        pl_gen34_redo_equalization;
  wire                        pl_gen34_redo_eq_speed;
  wire                        pl_gen34_eq_mismatch;



  wire [5:0]     pcie_rq_seq_num0_cc;
  wire           pcie_rq_seq_num_vld0_cc;

  // PCIE_4_0 Module
  generate
  if ((IMPL_TARGET == "SOFT") || (IMPL_TARGET == "PROTO")) begin  

  pcie_4_0_e4 #(

    .TCQ(TCQ)
   ,.IMPL_TARGET(IMPL_TARGET)
   ,.CRM_CORE_CLK_FREQ_500(CRM_CORE_CLK_FREQ_500)
   ,.CRM_USER_CLK_FREQ(CRM_USER_CLK_FREQ)
   ,.SIM_DEVICE(SIM_DEVICE)
   ,.AXISTEN_IF_WIDTH(AXISTEN_IF_WIDTH)
   ,.AXISTEN_IF_EXT_512(AXISTEN_IF_EXT_512)
   ,.AXISTEN_IF_EXT_512_CQ_STRADDLE(AXISTEN_IF_EXT_512_CQ_STRADDLE)
   ,.AXISTEN_IF_EXT_512_CC_STRADDLE(AXISTEN_IF_EXT_512_CC_STRADDLE)
   ,.AXISTEN_IF_EXT_512_RQ_STRADDLE(AXISTEN_IF_EXT_512_RQ_STRADDLE)
   ,.AXISTEN_IF_EXT_512_RC_STRADDLE(AXISTEN_IF_EXT_512_RC_STRADDLE)
   ,.AXISTEN_IF_CQ_ALIGNMENT_MODE(AXISTEN_IF_CQ_ALIGNMENT_MODE)
   ,.AXISTEN_IF_CC_ALIGNMENT_MODE(AXISTEN_IF_CC_ALIGNMENT_MODE)
   ,.AXISTEN_IF_RQ_ALIGNMENT_MODE(AXISTEN_IF_RQ_ALIGNMENT_MODE)
   ,.AXISTEN_IF_RC_ALIGNMENT_MODE(AXISTEN_IF_RC_ALIGNMENT_MODE)
   ,.AXISTEN_IF_RC_STRADDLE(AXISTEN_IF_RC_STRADDLE)
   ,.AXISTEN_IF_ENABLE_RX_MSG_INTFC(AXISTEN_IF_ENABLE_RX_MSG_INTFC)
   ,.AXISTEN_IF_ENABLE_MSG_ROUTE(AXISTEN_IF_ENABLE_MSG_ROUTE)
   ,.AXISTEN_IF_RX_PARITY_EN(AXISTEN_IF_RX_PARITY_EN)
   ,.AXISTEN_IF_TX_PARITY_EN(AXISTEN_IF_TX_PARITY_EN)
   ,.AXISTEN_IF_ENABLE_CLIENT_TAG(AXISTEN_IF_ENABLE_CLIENT_TAG)
   ,.AXISTEN_IF_ENABLE_256_TAGS(AXISTEN_IF_ENABLE_256_TAGS)
   ,.AXISTEN_IF_COMPL_TIMEOUT_REG0(AXISTEN_IF_COMPL_TIMEOUT_REG0)
   ,.AXISTEN_IF_COMPL_TIMEOUT_REG1(AXISTEN_IF_COMPL_TIMEOUT_REG1)
   ,.AXISTEN_IF_LEGACY_MODE_ENABLE(AXISTEN_IF_LEGACY_MODE_ENABLE)
   ,.AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK(AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK)
   ,.AXISTEN_IF_MSIX_TO_RAM_PIPELINE(AXISTEN_IF_MSIX_TO_RAM_PIPELINE)
   ,.AXISTEN_IF_MSIX_FROM_RAM_PIPELINE(AXISTEN_IF_MSIX_FROM_RAM_PIPELINE)
   ,.AXISTEN_IF_MSIX_RX_PARITY_EN(AXISTEN_IF_MSIX_RX_PARITY_EN)
   ,.AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE(AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE)
   ,.AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT(AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT)
   ,.AXISTEN_IF_CQ_EN_POISONED_MEM_WR(AXISTEN_IF_CQ_EN_POISONED_MEM_WR)
   ,.AXISTEN_IF_RQ_CC_REGISTERED_TREADY(AXISTEN_IF_RQ_CC_REGISTERED_TREADY)
   ,.PM_ASPML0S_TIMEOUT(PM_ASPML0S_TIMEOUT)
   ,.PM_L1_REENTRY_DELAY(PM_L1_REENTRY_DELAY)
   ,.PM_ASPML1_ENTRY_DELAY(PM_ASPML1_ENTRY_DELAY)
   ,.PM_ENABLE_SLOT_POWER_CAPTURE(PM_ENABLE_SLOT_POWER_CAPTURE)
   ,.PM_PME_SERVICE_TIMEOUT_DELAY(PM_PME_SERVICE_TIMEOUT_DELAY)
   ,.PM_PME_TURNOFF_ACK_DELAY(PM_PME_TURNOFF_ACK_DELAY)
   ,.PL_UPSTREAM_FACING(PL_UPSTREAM_FACING)
   ,.PL_LINK_CAP_MAX_LINK_WIDTH(PL_LINK_CAP_MAX_LINK_WIDTH)
   ,.PL_LINK_CAP_MAX_LINK_SPEED(PL_LINK_CAP_MAX_LINK_SPEED)
   ,.PL_DISABLE_DC_BALANCE(PL_DISABLE_DC_BALANCE)
   ,.PL_DISABLE_EI_INFER_IN_L0(PL_DISABLE_EI_INFER_IN_L0)
   ,.PL_N_FTS(PL_N_FTS)
   ,.PL_DISABLE_UPCONFIG_CAPABLE(PL_DISABLE_UPCONFIG_CAPABLE)
   ,.PL_DISABLE_RETRAIN_ON_FRAMING_ERROR(PL_DISABLE_RETRAIN_ON_FRAMING_ERROR)
   ,.PL_DISABLE_RETRAIN_ON_EB_ERROR(PL_DISABLE_RETRAIN_ON_EB_ERROR)
   ,.PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR(PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR)
   ,.PL_REPORT_ALL_PHY_ERRORS(PL_REPORT_ALL_PHY_ERRORS)
   ,.PL_DISABLE_LFSR_UPDATE_ON_SKP(PL_DISABLE_LFSR_UPDATE_ON_SKP)
   ,.PL_LANE0_EQ_CONTROL(PL_LANE0_EQ_CONTROL)
   ,.PL_LANE1_EQ_CONTROL(PL_LANE1_EQ_CONTROL)
   ,.PL_LANE2_EQ_CONTROL(PL_LANE2_EQ_CONTROL)
   ,.PL_LANE3_EQ_CONTROL(PL_LANE3_EQ_CONTROL)
   ,.PL_LANE4_EQ_CONTROL(PL_LANE4_EQ_CONTROL)
   ,.PL_LANE5_EQ_CONTROL(PL_LANE5_EQ_CONTROL)
   ,.PL_LANE6_EQ_CONTROL(PL_LANE6_EQ_CONTROL)
   ,.PL_LANE7_EQ_CONTROL(PL_LANE7_EQ_CONTROL)
   ,.PL_LANE8_EQ_CONTROL(PL_LANE8_EQ_CONTROL)
   ,.PL_LANE9_EQ_CONTROL(PL_LANE9_EQ_CONTROL)
   ,.PL_LANE10_EQ_CONTROL(PL_LANE10_EQ_CONTROL)
   ,.PL_LANE11_EQ_CONTROL(PL_LANE11_EQ_CONTROL)
   ,.PL_LANE12_EQ_CONTROL(PL_LANE12_EQ_CONTROL)
   ,.PL_LANE13_EQ_CONTROL(PL_LANE13_EQ_CONTROL)
   ,.PL_LANE14_EQ_CONTROL(PL_LANE14_EQ_CONTROL)
   ,.PL_LANE15_EQ_CONTROL(PL_LANE15_EQ_CONTROL)
   ,.PL_EQ_BYPASS_PHASE23(PL_EQ_BYPASS_PHASE23)
   ,.PL_EQ_ADAPT_ITER_COUNT(PL_EQ_ADAPT_ITER_COUNT)
   ,.PL_EQ_ADAPT_REJECT_RETRY_COUNT(PL_EQ_ADAPT_REJECT_RETRY_COUNT)
   ,.PL_EQ_SHORT_ADAPT_PHASE(PL_EQ_SHORT_ADAPT_PHASE)
   ,.PL_EQ_ADAPT_DISABLE_COEFF_CHECK(PL_EQ_ADAPT_DISABLE_COEFF_CHECK)
   ,.PL_EQ_ADAPT_DISABLE_PRESET_CHECK(PL_EQ_ADAPT_DISABLE_PRESET_CHECK)
   ,.PL_EQ_DEFAULT_TX_PRESET(PL_EQ_DEFAULT_TX_PRESET)
   ,.PL_EQ_DEFAULT_RX_PRESET_HINT(PL_EQ_DEFAULT_RX_PRESET_HINT)
   ,.PL_EQ_RX_ADAPT_EQ_PHASE0(PL_EQ_RX_ADAPT_EQ_PHASE0)
   ,.PL_EQ_RX_ADAPT_EQ_PHASE1(PL_EQ_RX_ADAPT_EQ_PHASE1)
   ,.PL_EQ_DISABLE_MISMATCH_CHECK(PL_EQ_DISABLE_MISMATCH_CHECK)
   ,.PL_RX_L0S_EXIT_TO_RECOVERY(PL_RX_L0S_EXIT_TO_RECOVERY)
   ,.PL_EQ_TX_8G_EQ_TS2_ENABLE(PL_EQ_TX_8G_EQ_TS2_ENABLE)
   ,.PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4(PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4)
   ,.PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3(PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3)
   ,.PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2(PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2)
   ,.PL_DESKEW_ON_SKIP_IN_GEN12(PL_DESKEW_ON_SKIP_IN_GEN12)
   ,.PL_INFER_EI_DISABLE_REC_RC(PL_INFER_EI_DISABLE_REC_RC)
   ,.PL_INFER_EI_DISABLE_REC_SPD(PL_INFER_EI_DISABLE_REC_SPD)
   ,.PL_INFER_EI_DISABLE_LPBK_ACTIVE(PL_INFER_EI_DISABLE_LPBK_ACTIVE)
   ,.PL_RX_ADAPT_TIMER_RRL_GEN3(PL_RX_ADAPT_TIMER_RRL_GEN3)
   ,.PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS(PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS)
   ,.PL_RX_ADAPT_TIMER_RRL_GEN4(PL_RX_ADAPT_TIMER_RRL_GEN4)
   ,.PL_RX_ADAPT_TIMER_CLWS_GEN3(PL_RX_ADAPT_TIMER_CLWS_GEN3)
   ,.PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS(PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS)
   ,.PL_RX_ADAPT_TIMER_CLWS_GEN4(PL_RX_ADAPT_TIMER_CLWS_GEN4)
   ,.PL_DISABLE_LANE_REVERSAL(PL_DISABLE_LANE_REVERSAL)
   ,.PL_CFG_STATE_ROBUSTNESS_ENABLE(PL_CFG_STATE_ROBUSTNESS_ENABLE)
   ,.PL_REDO_EQ_SOURCE_SELECT(PL_REDO_EQ_SOURCE_SELECT)
   ,.PL_DEEMPH_SOURCE_SELECT(PL_DEEMPH_SOURCE_SELECT)
   ,.PL_EXIT_LOOPBACK_ON_EI_ENTRY(PL_EXIT_LOOPBACK_ON_EI_ENTRY)
   ,.PL_QUIESCE_GUARANTEE_DISABLE(PL_QUIESCE_GUARANTEE_DISABLE)
   ,.PL_SRIS_ENABLE(PL_SRIS_ENABLE)
   ,.PL_SRIS_SKPOS_GEN_SPD_VEC(PL_SRIS_SKPOS_GEN_SPD_VEC)
   ,.PL_SRIS_SKPOS_REC_SPD_VEC(PL_SRIS_SKPOS_REC_SPD_VEC)
   ,.PL_SIM_FAST_LINK_TRAINING(PL_SIM_FAST_LINK_TRAINING)
   ,.PL_USER_SPARE(PL_USER_SPARE)
   ,.LL_ACK_TIMEOUT_EN(LL_ACK_TIMEOUT_EN)
   ,.LL_ACK_TIMEOUT(LL_ACK_TIMEOUT)
   ,.LL_ACK_TIMEOUT_FUNC(LL_ACK_TIMEOUT_FUNC)
   ,.LL_REPLAY_TIMEOUT_EN(LL_REPLAY_TIMEOUT_EN)
   ,.LL_REPLAY_TIMEOUT(LL_REPLAY_TIMEOUT)
   ,.LL_REPLAY_TIMEOUT_FUNC(LL_REPLAY_TIMEOUT_FUNC)
   ,.LL_REPLAY_TO_RAM_PIPELINE(LL_REPLAY_TO_RAM_PIPELINE)
   ,.LL_REPLAY_FROM_RAM_PIPELINE(LL_REPLAY_FROM_RAM_PIPELINE)
   ,.LL_DISABLE_SCHED_TX_NAK(LL_DISABLE_SCHED_TX_NAK)
   ,.LL_TX_TLP_PARITY_CHK(LL_TX_TLP_PARITY_CHK)
   ,.LL_RX_TLP_PARITY_GEN(LL_RX_TLP_PARITY_GEN)
   ,.LL_USER_SPARE(LL_USER_SPARE)
   ,.IS_SWITCH_PORT(IS_SWITCH_PORT)
   ,.CFG_BYPASS_MODE_ENABLE(CFG_BYPASS_MODE_ENABLE)
   ,.TL_PF_ENABLE_REG(TL_PF_ENABLE_REG)
   ,.TL_CREDITS_CD(TL_CREDITS_CD)
   ,.TL_CREDITS_CH(TL_CREDITS_CH)
   ,.TL_COMPLETION_RAM_SIZE(TL_COMPLETION_RAM_SIZE)
   ,.TL_COMPLETION_RAM_NUM_TLPS(TL_COMPLETION_RAM_NUM_TLPS)
   ,.TL_CREDITS_NPD(TL_CREDITS_NPD)
   ,.TL_CREDITS_NPH(TL_CREDITS_NPH)
   ,.TL_CREDITS_PD(TL_CREDITS_PD)
   ,.TL_CREDITS_PH(TL_CREDITS_PH)
   ,.TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE(TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE)
   ,.TL_RX_COMPLETION_TO_RAM_READ_PIPELINE(TL_RX_COMPLETION_TO_RAM_READ_PIPELINE)
   ,.TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE(TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE)
   ,.TL_POSTED_RAM_SIZE(TL_POSTED_RAM_SIZE)
   ,.TL_RX_POSTED_TO_RAM_WRITE_PIPELINE(TL_RX_POSTED_TO_RAM_WRITE_PIPELINE)
   ,.TL_RX_POSTED_TO_RAM_READ_PIPELINE(TL_RX_POSTED_TO_RAM_READ_PIPELINE)
   ,.TL_RX_POSTED_FROM_RAM_READ_PIPELINE(TL_RX_POSTED_FROM_RAM_READ_PIPELINE)
   ,.TL_TX_MUX_STRICT_PRIORITY(TL_TX_MUX_STRICT_PRIORITY)
   ,.TL_TX_TLP_STRADDLE_ENABLE(TL_TX_TLP_STRADDLE_ENABLE)
   ,.TL_TX_TLP_TERMINATE_PARITY(TL_TX_TLP_TERMINATE_PARITY)
   ,.TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT(TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT)
   ,.TL_FC_UPDATE_MIN_INTERVAL_TIME(TL_FC_UPDATE_MIN_INTERVAL_TIME)
   ,.TL_USER_SPARE(TL_USER_SPARE)
   ,.PF0_CLASS_CODE(PF0_CLASS_CODE)
   ,.PF1_CLASS_CODE(PF1_CLASS_CODE)
   ,.PF2_CLASS_CODE(PF2_CLASS_CODE)
   ,.PF3_CLASS_CODE(PF3_CLASS_CODE)
   ,.PF0_INTERRUPT_PIN(PF0_INTERRUPT_PIN)
   ,.PF1_INTERRUPT_PIN(PF1_INTERRUPT_PIN)
   ,.PF2_INTERRUPT_PIN(PF2_INTERRUPT_PIN)
   ,.PF3_INTERRUPT_PIN(PF3_INTERRUPT_PIN)
   ,.PF0_CAPABILITY_POINTER(PF0_CAPABILITY_POINTER)
   ,.PF1_CAPABILITY_POINTER(PF1_CAPABILITY_POINTER)
   ,.PF2_CAPABILITY_POINTER(PF2_CAPABILITY_POINTER)
   ,.PF3_CAPABILITY_POINTER(PF3_CAPABILITY_POINTER)
   ,.VF0_CAPABILITY_POINTER(VF0_CAPABILITY_POINTER)
   ,.LEGACY_CFG_EXTEND_INTERFACE_ENABLE(LEGACY_CFG_EXTEND_INTERFACE_ENABLE)
   ,.EXTENDED_CFG_EXTEND_INTERFACE_ENABLE(EXTENDED_CFG_EXTEND_INTERFACE_ENABLE)
   ,.TL2CFG_IF_PARITY_CHK(TL2CFG_IF_PARITY_CHK)
   ,.HEADER_TYPE_OVERRIDE(HEADER_TYPE_OVERRIDE)
   ,.PF0_BAR0_CONTROL(PF0_BAR0_CONTROL)
   ,.PF1_BAR0_CONTROL(PF1_BAR0_CONTROL)
   ,.PF2_BAR0_CONTROL(PF2_BAR0_CONTROL)
   ,.PF3_BAR0_CONTROL(PF3_BAR0_CONTROL)
   ,.PF0_BAR0_APERTURE_SIZE(PF0_BAR0_APERTURE_SIZE)
   ,.PF1_BAR0_APERTURE_SIZE(PF1_BAR0_APERTURE_SIZE)
   ,.PF2_BAR0_APERTURE_SIZE(PF2_BAR0_APERTURE_SIZE)
   ,.PF3_BAR0_APERTURE_SIZE(PF3_BAR0_APERTURE_SIZE)
   ,.PF0_BAR1_CONTROL(PF0_BAR1_CONTROL)
   ,.PF1_BAR1_CONTROL(PF1_BAR1_CONTROL)
   ,.PF2_BAR1_CONTROL(PF2_BAR1_CONTROL)
   ,.PF3_BAR1_CONTROL(PF3_BAR1_CONTROL)
   ,.PF0_BAR1_APERTURE_SIZE(PF0_BAR1_APERTURE_SIZE)
   ,.PF1_BAR1_APERTURE_SIZE(PF1_BAR1_APERTURE_SIZE)
   ,.PF2_BAR1_APERTURE_SIZE(PF2_BAR1_APERTURE_SIZE)
   ,.PF3_BAR1_APERTURE_SIZE(PF3_BAR1_APERTURE_SIZE)
   ,.PF0_BAR2_CONTROL(PF0_BAR2_CONTROL)
   ,.PF1_BAR2_CONTROL(PF1_BAR2_CONTROL)
   ,.PF2_BAR2_CONTROL(PF2_BAR2_CONTROL)
   ,.PF3_BAR2_CONTROL(PF3_BAR2_CONTROL)
   ,.PF0_BAR2_APERTURE_SIZE(PF0_BAR2_APERTURE_SIZE)
   ,.PF1_BAR2_APERTURE_SIZE(PF1_BAR2_APERTURE_SIZE)
   ,.PF2_BAR2_APERTURE_SIZE(PF2_BAR2_APERTURE_SIZE)
   ,.PF3_BAR2_APERTURE_SIZE(PF3_BAR2_APERTURE_SIZE)
   ,.PF0_BAR3_CONTROL(PF0_BAR3_CONTROL)
   ,.PF1_BAR3_CONTROL(PF1_BAR3_CONTROL)
   ,.PF2_BAR3_CONTROL(PF2_BAR3_CONTROL)
   ,.PF3_BAR3_CONTROL(PF3_BAR3_CONTROL)
   ,.PF0_BAR3_APERTURE_SIZE(PF0_BAR3_APERTURE_SIZE)
   ,.PF1_BAR3_APERTURE_SIZE(PF1_BAR3_APERTURE_SIZE)
   ,.PF2_BAR3_APERTURE_SIZE(PF2_BAR3_APERTURE_SIZE)
   ,.PF3_BAR3_APERTURE_SIZE(PF3_BAR3_APERTURE_SIZE)
   ,.PF0_BAR4_CONTROL(PF0_BAR4_CONTROL)
   ,.PF1_BAR4_CONTROL(PF1_BAR4_CONTROL)
   ,.PF2_BAR4_CONTROL(PF2_BAR4_CONTROL)
   ,.PF3_BAR4_CONTROL(PF3_BAR4_CONTROL)
   ,.PF0_BAR4_APERTURE_SIZE(PF0_BAR4_APERTURE_SIZE)
   ,.PF1_BAR4_APERTURE_SIZE(PF1_BAR4_APERTURE_SIZE)
   ,.PF2_BAR4_APERTURE_SIZE(PF2_BAR4_APERTURE_SIZE)
   ,.PF3_BAR4_APERTURE_SIZE(PF3_BAR4_APERTURE_SIZE)
   ,.PF0_BAR5_CONTROL(PF0_BAR5_CONTROL)
   ,.PF1_BAR5_CONTROL(PF1_BAR5_CONTROL)
   ,.PF2_BAR5_CONTROL(PF2_BAR5_CONTROL)
   ,.PF3_BAR5_CONTROL(PF3_BAR5_CONTROL)
   ,.PF0_BAR5_APERTURE_SIZE(PF0_BAR5_APERTURE_SIZE)
   ,.PF1_BAR5_APERTURE_SIZE(PF1_BAR5_APERTURE_SIZE)
   ,.PF2_BAR5_APERTURE_SIZE(PF2_BAR5_APERTURE_SIZE)
   ,.PF3_BAR5_APERTURE_SIZE(PF3_BAR5_APERTURE_SIZE)
   ,.PF0_EXPANSION_ROM_ENABLE(PF0_EXPANSION_ROM_ENABLE)
   ,.PF1_EXPANSION_ROM_ENABLE(PF1_EXPANSION_ROM_ENABLE)
   ,.PF2_EXPANSION_ROM_ENABLE(PF2_EXPANSION_ROM_ENABLE)
   ,.PF3_EXPANSION_ROM_ENABLE(PF3_EXPANSION_ROM_ENABLE)
   ,.PF0_EXPANSION_ROM_APERTURE_SIZE(PF0_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF1_EXPANSION_ROM_APERTURE_SIZE(PF1_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF2_EXPANSION_ROM_APERTURE_SIZE(PF2_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF3_EXPANSION_ROM_APERTURE_SIZE(PF3_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF0_PCIE_CAP_NEXTPTR(PF0_PCIE_CAP_NEXTPTR)
   ,.PF1_PCIE_CAP_NEXTPTR(PF1_PCIE_CAP_NEXTPTR)
   ,.PF2_PCIE_CAP_NEXTPTR(PF2_PCIE_CAP_NEXTPTR)
   ,.PF3_PCIE_CAP_NEXTPTR(PF3_PCIE_CAP_NEXTPTR)
   ,.VFG0_PCIE_CAP_NEXTPTR(VFG0_PCIE_CAP_NEXTPTR)
   ,.VFG1_PCIE_CAP_NEXTPTR(VFG1_PCIE_CAP_NEXTPTR)
   ,.VFG2_PCIE_CAP_NEXTPTR(VFG2_PCIE_CAP_NEXTPTR)
   ,.VFG3_PCIE_CAP_NEXTPTR(VFG3_PCIE_CAP_NEXTPTR)
   ,.PF0_DEV_CAP_MAX_PAYLOAD_SIZE(PF0_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF1_DEV_CAP_MAX_PAYLOAD_SIZE(PF1_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF2_DEV_CAP_MAX_PAYLOAD_SIZE(PF2_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF3_DEV_CAP_MAX_PAYLOAD_SIZE(PF3_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF0_DEV_CAP_EXT_TAG_SUPPORTED(PF0_DEV_CAP_EXT_TAG_SUPPORTED)
   ,.PF0_DEV_CAP_ENDPOINT_L0S_LATENCY(PF0_DEV_CAP_ENDPOINT_L0S_LATENCY)
   ,.PF0_DEV_CAP_ENDPOINT_L1_LATENCY(PF0_DEV_CAP_ENDPOINT_L1_LATENCY)
   ,.PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE(PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE)
   ,.PF0_LINK_CAP_ASPM_SUPPORT(PF0_LINK_CAP_ASPM_SUPPORT)
   ,.PF0_LINK_CONTROL_RCB(PF0_LINK_CONTROL_RCB)
   ,.PF0_LINK_STATUS_SLOT_CLOCK_CONFIG(PF0_LINK_STATUS_SLOT_CLOCK_CONFIG)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4)
   ,.PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE(PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE)
   ,.PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT(PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT(PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT(PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_LTR_SUPPORT(PF0_DEV_CAP2_LTR_SUPPORT)
   ,.PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT(PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_OBFF_SUPPORT(PF0_DEV_CAP2_OBFF_SUPPORT)
   ,.PF0_DEV_CAP2_ARI_FORWARD_ENABLE(PF0_DEV_CAP2_ARI_FORWARD_ENABLE)
   ,.PF0_MSI_CAP_NEXTPTR(PF0_MSI_CAP_NEXTPTR)
   ,.PF1_MSI_CAP_NEXTPTR(PF1_MSI_CAP_NEXTPTR)
   ,.PF2_MSI_CAP_NEXTPTR(PF2_MSI_CAP_NEXTPTR)
   ,.PF3_MSI_CAP_NEXTPTR(PF3_MSI_CAP_NEXTPTR)
   ,.PF0_MSI_CAP_PERVECMASKCAP(PF0_MSI_CAP_PERVECMASKCAP)
   ,.PF1_MSI_CAP_PERVECMASKCAP(PF1_MSI_CAP_PERVECMASKCAP)
   ,.PF2_MSI_CAP_PERVECMASKCAP(PF2_MSI_CAP_PERVECMASKCAP)
   ,.PF3_MSI_CAP_PERVECMASKCAP(PF3_MSI_CAP_PERVECMASKCAP)
   ,.PF0_MSI_CAP_MULTIMSGCAP(PF0_MSI_CAP_MULTIMSGCAP)
   ,.PF1_MSI_CAP_MULTIMSGCAP(PF1_MSI_CAP_MULTIMSGCAP)
   ,.PF2_MSI_CAP_MULTIMSGCAP(PF2_MSI_CAP_MULTIMSGCAP)
   ,.PF3_MSI_CAP_MULTIMSGCAP(PF3_MSI_CAP_MULTIMSGCAP)
   ,.PF0_MSIX_CAP_NEXTPTR(PF0_MSIX_CAP_NEXTPTR)
   ,.PF1_MSIX_CAP_NEXTPTR(PF1_MSIX_CAP_NEXTPTR)
   ,.PF2_MSIX_CAP_NEXTPTR(PF2_MSIX_CAP_NEXTPTR)
   ,.PF3_MSIX_CAP_NEXTPTR(PF3_MSIX_CAP_NEXTPTR)
   ,.VFG0_MSIX_CAP_NEXTPTR(VFG0_MSIX_CAP_NEXTPTR)
   ,.VFG1_MSIX_CAP_NEXTPTR(VFG1_MSIX_CAP_NEXTPTR)
   ,.VFG2_MSIX_CAP_NEXTPTR(VFG2_MSIX_CAP_NEXTPTR)
   ,.VFG3_MSIX_CAP_NEXTPTR(VFG3_MSIX_CAP_NEXTPTR)
   ,.PF0_MSIX_CAP_PBA_BIR(PF0_MSIX_CAP_PBA_BIR)
   ,.PF1_MSIX_CAP_PBA_BIR(PF1_MSIX_CAP_PBA_BIR)
   ,.PF2_MSIX_CAP_PBA_BIR(PF2_MSIX_CAP_PBA_BIR)
   ,.PF3_MSIX_CAP_PBA_BIR(PF3_MSIX_CAP_PBA_BIR)
   ,.VFG0_MSIX_CAP_PBA_BIR(VFG0_MSIX_CAP_PBA_BIR)
   ,.VFG1_MSIX_CAP_PBA_BIR(VFG1_MSIX_CAP_PBA_BIR)
   ,.VFG2_MSIX_CAP_PBA_BIR(VFG2_MSIX_CAP_PBA_BIR)
   ,.VFG3_MSIX_CAP_PBA_BIR(VFG3_MSIX_CAP_PBA_BIR)
   ,.PF0_MSIX_CAP_PBA_OFFSET(PF0_MSIX_CAP_PBA_OFFSET)
   ,.PF1_MSIX_CAP_PBA_OFFSET(PF1_MSIX_CAP_PBA_OFFSET)
   ,.PF2_MSIX_CAP_PBA_OFFSET(PF2_MSIX_CAP_PBA_OFFSET)
   ,.PF3_MSIX_CAP_PBA_OFFSET(PF3_MSIX_CAP_PBA_OFFSET)
   ,.VFG0_MSIX_CAP_PBA_OFFSET(VFG0_MSIX_CAP_PBA_OFFSET)
   ,.VFG1_MSIX_CAP_PBA_OFFSET(VFG1_MSIX_CAP_PBA_OFFSET)
   ,.VFG2_MSIX_CAP_PBA_OFFSET(VFG2_MSIX_CAP_PBA_OFFSET)
   ,.VFG3_MSIX_CAP_PBA_OFFSET(VFG3_MSIX_CAP_PBA_OFFSET)
   ,.PF0_MSIX_CAP_TABLE_BIR(PF0_MSIX_CAP_TABLE_BIR)
   ,.PF1_MSIX_CAP_TABLE_BIR(PF1_MSIX_CAP_TABLE_BIR)
   ,.PF2_MSIX_CAP_TABLE_BIR(PF2_MSIX_CAP_TABLE_BIR)
   ,.PF3_MSIX_CAP_TABLE_BIR(PF3_MSIX_CAP_TABLE_BIR)
   ,.VFG0_MSIX_CAP_TABLE_BIR(VFG0_MSIX_CAP_TABLE_BIR)
   ,.VFG1_MSIX_CAP_TABLE_BIR(VFG1_MSIX_CAP_TABLE_BIR)
   ,.VFG2_MSIX_CAP_TABLE_BIR(VFG2_MSIX_CAP_TABLE_BIR)
   ,.VFG3_MSIX_CAP_TABLE_BIR(VFG3_MSIX_CAP_TABLE_BIR)
   ,.PF0_MSIX_CAP_TABLE_OFFSET(PF0_MSIX_CAP_TABLE_OFFSET)
   ,.PF1_MSIX_CAP_TABLE_OFFSET(PF1_MSIX_CAP_TABLE_OFFSET)
   ,.PF2_MSIX_CAP_TABLE_OFFSET(PF2_MSIX_CAP_TABLE_OFFSET)
   ,.PF3_MSIX_CAP_TABLE_OFFSET(PF3_MSIX_CAP_TABLE_OFFSET)
   ,.VFG0_MSIX_CAP_TABLE_OFFSET(VFG0_MSIX_CAP_TABLE_OFFSET)
   ,.VFG1_MSIX_CAP_TABLE_OFFSET(VFG1_MSIX_CAP_TABLE_OFFSET)
   ,.VFG2_MSIX_CAP_TABLE_OFFSET(VFG2_MSIX_CAP_TABLE_OFFSET)
   ,.VFG3_MSIX_CAP_TABLE_OFFSET(VFG3_MSIX_CAP_TABLE_OFFSET)
   ,.PF0_MSIX_CAP_TABLE_SIZE(PF0_MSIX_CAP_TABLE_SIZE)
   ,.PF1_MSIX_CAP_TABLE_SIZE(PF1_MSIX_CAP_TABLE_SIZE)
   ,.PF2_MSIX_CAP_TABLE_SIZE(PF2_MSIX_CAP_TABLE_SIZE)
   ,.PF3_MSIX_CAP_TABLE_SIZE(PF3_MSIX_CAP_TABLE_SIZE)
   ,.VFG0_MSIX_CAP_TABLE_SIZE(VFG0_MSIX_CAP_TABLE_SIZE)
   ,.VFG1_MSIX_CAP_TABLE_SIZE(VFG1_MSIX_CAP_TABLE_SIZE)
   ,.VFG2_MSIX_CAP_TABLE_SIZE(VFG2_MSIX_CAP_TABLE_SIZE)
   ,.VFG3_MSIX_CAP_TABLE_SIZE(VFG3_MSIX_CAP_TABLE_SIZE)
   ,.PF0_MSIX_VECTOR_COUNT(PF0_MSIX_VECTOR_COUNT)
   ,.PF0_PM_CAP_ID(PF0_PM_CAP_ID)
   ,.PF0_PM_CAP_NEXTPTR(PF0_PM_CAP_NEXTPTR)
   ,.PF1_PM_CAP_NEXTPTR(PF1_PM_CAP_NEXTPTR)
   ,.PF2_PM_CAP_NEXTPTR(PF2_PM_CAP_NEXTPTR)
   ,.PF3_PM_CAP_NEXTPTR(PF3_PM_CAP_NEXTPTR)
   ,.PF0_PM_CAP_PMESUPPORT_D3HOT(PF0_PM_CAP_PMESUPPORT_D3HOT)
   ,.PF0_PM_CAP_PMESUPPORT_D1(PF0_PM_CAP_PMESUPPORT_D1)
   ,.PF0_PM_CAP_PMESUPPORT_D0(PF0_PM_CAP_PMESUPPORT_D0)
   ,.PF0_PM_CAP_SUPP_D1_STATE(PF0_PM_CAP_SUPP_D1_STATE)
   ,.PF0_PM_CAP_VER_ID(PF0_PM_CAP_VER_ID)
   ,.PF0_PM_CSR_NOSOFTRESET(PF0_PM_CSR_NOSOFTRESET)
   ,.PM_ENABLE_L23_ENTRY(PM_ENABLE_L23_ENTRY)
   ,.DNSTREAM_LINK_NUM(DNSTREAM_LINK_NUM)
   ,.AUTO_FLR_RESPONSE(AUTO_FLR_RESPONSE)
   ,.PF0_DSN_CAP_NEXTPTR(PF0_DSN_CAP_NEXTPTR)
   ,.PF1_DSN_CAP_NEXTPTR(PF1_DSN_CAP_NEXTPTR)
   ,.PF2_DSN_CAP_NEXTPTR(PF2_DSN_CAP_NEXTPTR)
   ,.PF3_DSN_CAP_NEXTPTR(PF3_DSN_CAP_NEXTPTR)
   ,.DSN_CAP_ENABLE(DSN_CAP_ENABLE)
   ,.PF0_VC_CAP_VER(PF0_VC_CAP_VER)
   ,.PF0_VC_CAP_NEXTPTR(PF0_VC_CAP_NEXTPTR)
   ,.PF0_VC_CAP_ENABLE(PF0_VC_CAP_ENABLE)
   ,.PF0_SECONDARY_PCIE_CAP_NEXTPTR(PF0_SECONDARY_PCIE_CAP_NEXTPTR)
   ,.PF0_AER_CAP_NEXTPTR(PF0_AER_CAP_NEXTPTR)
   ,.PF1_AER_CAP_NEXTPTR(PF1_AER_CAP_NEXTPTR)
   ,.PF2_AER_CAP_NEXTPTR(PF2_AER_CAP_NEXTPTR)
   ,.PF3_AER_CAP_NEXTPTR(PF3_AER_CAP_NEXTPTR)
   ,.PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE(PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE)
   ,.ARI_CAP_ENABLE(ARI_CAP_ENABLE)
   ,.PF0_ARI_CAP_NEXTPTR(PF0_ARI_CAP_NEXTPTR)
   ,.PF1_ARI_CAP_NEXTPTR(PF1_ARI_CAP_NEXTPTR)
   ,.PF2_ARI_CAP_NEXTPTR(PF2_ARI_CAP_NEXTPTR)
   ,.PF3_ARI_CAP_NEXTPTR(PF3_ARI_CAP_NEXTPTR)
   ,.VFG0_ARI_CAP_NEXTPTR(VFG0_ARI_CAP_NEXTPTR)
   ,.VFG1_ARI_CAP_NEXTPTR(VFG1_ARI_CAP_NEXTPTR)
   ,.VFG2_ARI_CAP_NEXTPTR(VFG2_ARI_CAP_NEXTPTR)
   ,.VFG3_ARI_CAP_NEXTPTR(VFG3_ARI_CAP_NEXTPTR)
   ,.PF0_ARI_CAP_VER(PF0_ARI_CAP_VER)
   ,.PF0_ARI_CAP_NEXT_FUNC(PF0_ARI_CAP_NEXT_FUNC)
   ,.PF1_ARI_CAP_NEXT_FUNC(PF1_ARI_CAP_NEXT_FUNC)
   ,.PF2_ARI_CAP_NEXT_FUNC(PF2_ARI_CAP_NEXT_FUNC)
   ,.PF3_ARI_CAP_NEXT_FUNC(PF3_ARI_CAP_NEXT_FUNC)
   ,.PF0_LTR_CAP_NEXTPTR(PF0_LTR_CAP_NEXTPTR)
   ,.PF0_LTR_CAP_VER(PF0_LTR_CAP_VER)
   ,.PF0_LTR_CAP_MAX_SNOOP_LAT(PF0_LTR_CAP_MAX_SNOOP_LAT)
   ,.PF0_LTR_CAP_MAX_NOSNOOP_LAT(PF0_LTR_CAP_MAX_NOSNOOP_LAT)
   ,.LTR_TX_MESSAGE_ON_LTR_ENABLE(LTR_TX_MESSAGE_ON_LTR_ENABLE)
   ,.LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE(LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE)
   ,.LTR_TX_MESSAGE_MINIMUM_INTERVAL(LTR_TX_MESSAGE_MINIMUM_INTERVAL)
   ,.SRIOV_CAP_ENABLE(SRIOV_CAP_ENABLE)
   ,.PF0_SRIOV_CAP_NEXTPTR(PF0_SRIOV_CAP_NEXTPTR)
   ,.PF1_SRIOV_CAP_NEXTPTR(PF1_SRIOV_CAP_NEXTPTR)
   ,.PF2_SRIOV_CAP_NEXTPTR(PF2_SRIOV_CAP_NEXTPTR)
   ,.PF3_SRIOV_CAP_NEXTPTR(PF3_SRIOV_CAP_NEXTPTR)
   ,.PF0_SRIOV_CAP_VER(PF0_SRIOV_CAP_VER)
   ,.PF1_SRIOV_CAP_VER(PF1_SRIOV_CAP_VER)
   ,.PF2_SRIOV_CAP_VER(PF2_SRIOV_CAP_VER)
   ,.PF3_SRIOV_CAP_VER(PF3_SRIOV_CAP_VER)
   ,.PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF0_SRIOV_CAP_INITIAL_VF(PF0_SRIOV_CAP_INITIAL_VF)
   ,.PF1_SRIOV_CAP_INITIAL_VF(PF1_SRIOV_CAP_INITIAL_VF)
   ,.PF2_SRIOV_CAP_INITIAL_VF(PF2_SRIOV_CAP_INITIAL_VF)
   ,.PF3_SRIOV_CAP_INITIAL_VF(PF3_SRIOV_CAP_INITIAL_VF)
   ,.PF0_SRIOV_CAP_TOTAL_VF(PF0_SRIOV_CAP_TOTAL_VF)
   ,.PF1_SRIOV_CAP_TOTAL_VF(PF1_SRIOV_CAP_TOTAL_VF)
   ,.PF2_SRIOV_CAP_TOTAL_VF(PF2_SRIOV_CAP_TOTAL_VF)
   ,.PF3_SRIOV_CAP_TOTAL_VF(PF3_SRIOV_CAP_TOTAL_VF)
   ,.PF0_SRIOV_FUNC_DEP_LINK(PF0_SRIOV_FUNC_DEP_LINK)
   ,.PF1_SRIOV_FUNC_DEP_LINK(PF1_SRIOV_FUNC_DEP_LINK)
   ,.PF2_SRIOV_FUNC_DEP_LINK(PF2_SRIOV_FUNC_DEP_LINK)
   ,.PF3_SRIOV_FUNC_DEP_LINK(PF3_SRIOV_FUNC_DEP_LINK)
   ,.PF0_SRIOV_FIRST_VF_OFFSET(PF0_SRIOV_FIRST_VF_OFFSET)
   ,.PF1_SRIOV_FIRST_VF_OFFSET(PF1_SRIOV_FIRST_VF_OFFSET)
   ,.PF2_SRIOV_FIRST_VF_OFFSET(PF2_SRIOV_FIRST_VF_OFFSET)
   ,.PF3_SRIOV_FIRST_VF_OFFSET(PF3_SRIOV_FIRST_VF_OFFSET)
   ,.PF0_SRIOV_VF_DEVICE_ID(PF0_SRIOV_VF_DEVICE_ID)
   ,.PF1_SRIOV_VF_DEVICE_ID(PF1_SRIOV_VF_DEVICE_ID)
   ,.PF2_SRIOV_VF_DEVICE_ID(PF2_SRIOV_VF_DEVICE_ID)
   ,.PF3_SRIOV_VF_DEVICE_ID(PF3_SRIOV_VF_DEVICE_ID)
   ,.PF0_SRIOV_SUPPORTED_PAGE_SIZE(PF0_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF1_SRIOV_SUPPORTED_PAGE_SIZE(PF1_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF2_SRIOV_SUPPORTED_PAGE_SIZE(PF2_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF3_SRIOV_SUPPORTED_PAGE_SIZE(PF3_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF0_SRIOV_BAR0_CONTROL(PF0_SRIOV_BAR0_CONTROL)
   ,.PF1_SRIOV_BAR0_CONTROL(PF1_SRIOV_BAR0_CONTROL)
   ,.PF2_SRIOV_BAR0_CONTROL(PF2_SRIOV_BAR0_CONTROL)
   ,.PF3_SRIOV_BAR0_CONTROL(PF3_SRIOV_BAR0_CONTROL)
   ,.PF0_SRIOV_BAR0_APERTURE_SIZE(PF0_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR0_APERTURE_SIZE(PF1_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR0_APERTURE_SIZE(PF2_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR0_APERTURE_SIZE(PF3_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR1_CONTROL(PF0_SRIOV_BAR1_CONTROL)
   ,.PF1_SRIOV_BAR1_CONTROL(PF1_SRIOV_BAR1_CONTROL)
   ,.PF2_SRIOV_BAR1_CONTROL(PF2_SRIOV_BAR1_CONTROL)
   ,.PF3_SRIOV_BAR1_CONTROL(PF3_SRIOV_BAR1_CONTROL)
   ,.PF0_SRIOV_BAR1_APERTURE_SIZE(PF0_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR1_APERTURE_SIZE(PF1_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR1_APERTURE_SIZE(PF2_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR1_APERTURE_SIZE(PF3_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR2_CONTROL(PF0_SRIOV_BAR2_CONTROL)
   ,.PF1_SRIOV_BAR2_CONTROL(PF1_SRIOV_BAR2_CONTROL)
   ,.PF2_SRIOV_BAR2_CONTROL(PF2_SRIOV_BAR2_CONTROL)
   ,.PF3_SRIOV_BAR2_CONTROL(PF3_SRIOV_BAR2_CONTROL)
   ,.PF0_SRIOV_BAR2_APERTURE_SIZE(PF0_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR2_APERTURE_SIZE(PF1_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR2_APERTURE_SIZE(PF2_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR2_APERTURE_SIZE(PF3_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR3_CONTROL(PF0_SRIOV_BAR3_CONTROL)
   ,.PF1_SRIOV_BAR3_CONTROL(PF1_SRIOV_BAR3_CONTROL)
   ,.PF2_SRIOV_BAR3_CONTROL(PF2_SRIOV_BAR3_CONTROL)
   ,.PF3_SRIOV_BAR3_CONTROL(PF3_SRIOV_BAR3_CONTROL)
   ,.PF0_SRIOV_BAR3_APERTURE_SIZE(PF0_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR3_APERTURE_SIZE(PF1_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR3_APERTURE_SIZE(PF2_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR3_APERTURE_SIZE(PF3_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR4_CONTROL(PF0_SRIOV_BAR4_CONTROL)
   ,.PF1_SRIOV_BAR4_CONTROL(PF1_SRIOV_BAR4_CONTROL)
   ,.PF2_SRIOV_BAR4_CONTROL(PF2_SRIOV_BAR4_CONTROL)
   ,.PF3_SRIOV_BAR4_CONTROL(PF3_SRIOV_BAR4_CONTROL)
   ,.PF0_SRIOV_BAR4_APERTURE_SIZE(PF0_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR4_APERTURE_SIZE(PF1_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR4_APERTURE_SIZE(PF2_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR4_APERTURE_SIZE(PF3_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR5_CONTROL(PF0_SRIOV_BAR5_CONTROL)
   ,.PF1_SRIOV_BAR5_CONTROL(PF1_SRIOV_BAR5_CONTROL)
   ,.PF2_SRIOV_BAR5_CONTROL(PF2_SRIOV_BAR5_CONTROL)
   ,.PF3_SRIOV_BAR5_CONTROL(PF3_SRIOV_BAR5_CONTROL)
   ,.PF0_SRIOV_BAR5_APERTURE_SIZE(PF0_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR5_APERTURE_SIZE(PF1_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR5_APERTURE_SIZE(PF2_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR5_APERTURE_SIZE(PF3_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF0_TPHR_CAP_NEXTPTR(PF0_TPHR_CAP_NEXTPTR)
   ,.PF1_TPHR_CAP_NEXTPTR(PF1_TPHR_CAP_NEXTPTR)
   ,.PF2_TPHR_CAP_NEXTPTR(PF2_TPHR_CAP_NEXTPTR)
   ,.PF3_TPHR_CAP_NEXTPTR(PF3_TPHR_CAP_NEXTPTR)
   ,.VFG0_TPHR_CAP_NEXTPTR(VFG0_TPHR_CAP_NEXTPTR)
   ,.VFG1_TPHR_CAP_NEXTPTR(VFG1_TPHR_CAP_NEXTPTR)
   ,.VFG2_TPHR_CAP_NEXTPTR(VFG2_TPHR_CAP_NEXTPTR)
   ,.VFG3_TPHR_CAP_NEXTPTR(VFG3_TPHR_CAP_NEXTPTR)
   ,.PF0_TPHR_CAP_VER(PF0_TPHR_CAP_VER)
   ,.PF0_TPHR_CAP_INT_VEC_MODE(PF0_TPHR_CAP_INT_VEC_MODE)
   ,.PF0_TPHR_CAP_DEV_SPECIFIC_MODE(PF0_TPHR_CAP_DEV_SPECIFIC_MODE)
   ,.PF0_TPHR_CAP_ST_TABLE_LOC(PF0_TPHR_CAP_ST_TABLE_LOC)
   ,.PF0_TPHR_CAP_ST_TABLE_SIZE(PF0_TPHR_CAP_ST_TABLE_SIZE)
   ,.PF0_TPHR_CAP_ST_MODE_SEL(PF0_TPHR_CAP_ST_MODE_SEL)
   ,.PF1_TPHR_CAP_ST_MODE_SEL(PF1_TPHR_CAP_ST_MODE_SEL)
   ,.PF2_TPHR_CAP_ST_MODE_SEL(PF2_TPHR_CAP_ST_MODE_SEL)
   ,.PF3_TPHR_CAP_ST_MODE_SEL(PF3_TPHR_CAP_ST_MODE_SEL)
   ,.VFG0_TPHR_CAP_ST_MODE_SEL(VFG0_TPHR_CAP_ST_MODE_SEL)
   ,.VFG1_TPHR_CAP_ST_MODE_SEL(VFG1_TPHR_CAP_ST_MODE_SEL)
   ,.VFG2_TPHR_CAP_ST_MODE_SEL(VFG2_TPHR_CAP_ST_MODE_SEL)
   ,.VFG3_TPHR_CAP_ST_MODE_SEL(VFG3_TPHR_CAP_ST_MODE_SEL)
   ,.PF0_TPHR_CAP_ENABLE(PF0_TPHR_CAP_ENABLE)
   ,.TPH_TO_RAM_PIPELINE(TPH_TO_RAM_PIPELINE)
   ,.TPH_FROM_RAM_PIPELINE(TPH_FROM_RAM_PIPELINE)
   ,.MCAP_ENABLE(MCAP_ENABLE)
   ,.MCAP_CONFIGURE_OVERRIDE(MCAP_CONFIGURE_OVERRIDE)
   ,.MCAP_CAP_NEXTPTR(MCAP_CAP_NEXTPTR)
   ,.MCAP_VSEC_ID(MCAP_VSEC_ID)
   ,.MCAP_VSEC_REV(MCAP_VSEC_REV)
   ,.MCAP_VSEC_LEN(MCAP_VSEC_LEN)
   ,.MCAP_FPGA_BITSTREAM_VERSION(MCAP_FPGA_BITSTREAM_VERSION)
   ,.MCAP_INTERRUPT_ON_MCAP_EOS(MCAP_INTERRUPT_ON_MCAP_EOS)
   ,.MCAP_INTERRUPT_ON_MCAP_ERROR(MCAP_INTERRUPT_ON_MCAP_ERROR)
   ,.MCAP_INPUT_GATE_DESIGN_SWITCH(MCAP_INPUT_GATE_DESIGN_SWITCH)
   ,.MCAP_EOS_DESIGN_SWITCH(MCAP_EOS_DESIGN_SWITCH)
   ,.MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH(MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH)
   ,.MCAP_GATE_IO_ENABLE_DESIGN_SWITCH(MCAP_GATE_IO_ENABLE_DESIGN_SWITCH)
   ,.SIM_JTAG_IDCODE(SIM_JTAG_IDCODE)
   ,.DEBUG_AXIST_DISABLE_FEATURE_BIT(DEBUG_AXIST_DISABLE_FEATURE_BIT)
   ,.DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS(DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS)
   ,.DEBUG_TL_DISABLE_FC_TIMEOUT(DEBUG_TL_DISABLE_FC_TIMEOUT)
   ,.DEBUG_PL_DISABLE_SCRAMBLING(DEBUG_PL_DISABLE_SCRAMBLING)
   ,.DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL (DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL )
   ,.DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW (DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW )
   ,.DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR(DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR)
   ,.DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR(DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR)
   ,.DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR(DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR)
   ,.DEBUG_PL_SIM_RESET_LFSR(DEBUG_PL_SIM_RESET_LFSR)
   ,.DEBUG_PL_SPARE(DEBUG_PL_SPARE)
   ,.DEBUG_LL_SPARE(DEBUG_LL_SPARE)
   ,.DEBUG_TL_SPARE(DEBUG_TL_SPARE)
   ,.DEBUG_AXI4ST_SPARE(DEBUG_AXI4ST_SPARE)
   ,.DEBUG_CFG_SPARE(DEBUG_CFG_SPARE)
   ,.DEBUG_CAR_SPARE(DEBUG_CAR_SPARE)
   ,.TEST_MODE_PIN_CHAR(TEST_MODE_PIN_CHAR)
   ,.SPARE_BIT0(SPARE_BIT0)
   ,.SPARE_BIT1(SPARE_BIT1)
   ,.SPARE_BIT2(SPARE_BIT2)
   ,.SPARE_BIT3(SPARE_BIT3)
   ,.SPARE_BIT4(SPARE_BIT4)
   ,.SPARE_BIT5(SPARE_BIT5)
   ,.SPARE_BIT6(SPARE_BIT6)
   ,.SPARE_BIT7(SPARE_BIT7)
   ,.SPARE_BIT8(SPARE_BIT8)
   ,.SPARE_BYTE0(SPARE_BYTE0)
   ,.SPARE_BYTE1(SPARE_BYTE1)
   ,.SPARE_BYTE2(SPARE_BYTE2)
   ,.SPARE_BYTE3(SPARE_BYTE3)
   ,.SPARE_WORD0(SPARE_WORD0)
   ,.SPARE_WORD1(SPARE_WORD1)
   ,.SPARE_WORD2(SPARE_WORD2)
   ,.SPARE_WORD3(SPARE_WORD3)

  ) pcie_4_0_e4_inst ( 

    .mi_replay_ram_address0(mi_replay_ram_address0[8:0])
   ,.mi_replay_ram_address1(mi_replay_ram_address1[8:0])
   ,.mi_replay_ram_write_data0(mi_replay_ram_write_data0[127:0])
   ,.mi_replay_ram_write_enable0(mi_replay_ram_write_enable0)
   ,.mi_replay_ram_write_data1(mi_replay_ram_write_data1[127:0])
   ,.mi_replay_ram_write_enable1(mi_replay_ram_write_enable1)
   ,.mi_replay_ram_read_data0(mi_replay_ram_read_data0[127:0])
   ,.mi_replay_ram_read_enable0(mi_replay_ram_read_enable0)
   ,.mi_replay_ram_read_data1(mi_replay_ram_read_data1[127:0])
   ,.mi_replay_ram_read_enable1(mi_replay_ram_read_enable1)
   ,.mi_replay_ram_err_cor(mi_replay_ram_err_cor[5:0])
   ,.mi_replay_ram_err_uncor(mi_replay_ram_err_uncor[5:0])
   ,.mi_rx_posted_request_ram_write_address0(mi_rx_posted_request_ram_write_address0[8:0])
   ,.mi_rx_posted_request_ram_write_data0(mi_rx_posted_request_ram_write_data0[143:0])
   ,.mi_rx_posted_request_ram_write_enable0(mi_rx_posted_request_ram_write_enable0)
   ,.mi_rx_posted_request_ram_write_address1(mi_rx_posted_request_ram_write_address1[8:0])
   ,.mi_rx_posted_request_ram_write_data1(mi_rx_posted_request_ram_write_data1[143:0])
   ,.mi_rx_posted_request_ram_write_enable1(mi_rx_posted_request_ram_write_enable1)
   ,.mi_rx_posted_request_ram_read_address0(mi_rx_posted_request_ram_read_address0[8:0])
   ,.mi_rx_posted_request_ram_read_data0(mi_rx_posted_request_ram_read_data0[143:0])
   ,.mi_rx_posted_request_ram_read_enable0(mi_rx_posted_request_ram_read_enable0)
   ,.mi_rx_posted_request_ram_read_address1(mi_rx_posted_request_ram_read_address1[8:0])
   ,.mi_rx_posted_request_ram_read_data1(mi_rx_posted_request_ram_read_data1[143:0])
   ,.mi_rx_posted_request_ram_read_enable1(mi_rx_posted_request_ram_read_enable1)
   ,.mi_rx_posted_request_ram_err_cor(mi_rx_posted_request_ram_err_cor[5:0])
   ,.mi_rx_posted_request_ram_err_uncor(mi_rx_posted_request_ram_err_uncor[5:0])
   ,.mi_rx_completion_ram_write_address0(mi_rx_completion_ram_write_address0[8:0])
   ,.mi_rx_completion_ram_write_data0(mi_rx_completion_ram_write_data0[143:0])
   ,.mi_rx_completion_ram_write_enable0(mi_rx_completion_ram_write_enable0[1:0])
   ,.mi_rx_completion_ram_write_address1(mi_rx_completion_ram_write_address1[8:0])
   ,.mi_rx_completion_ram_write_data1(mi_rx_completion_ram_write_data1[143:0])
   ,.mi_rx_completion_ram_write_enable1(mi_rx_completion_ram_write_enable1[1:0])
   ,.mi_rx_completion_ram_read_address0(mi_rx_completion_ram_read_address0[8:0])
   ,.mi_rx_completion_ram_read_data0(mi_rx_completion_ram_read_data0[143:0])
   ,.mi_rx_completion_ram_read_enable0(mi_rx_completion_ram_read_enable0[1:0])
   ,.mi_rx_completion_ram_read_address1(mi_rx_completion_ram_read_address1[8:0])
   ,.mi_rx_completion_ram_read_data1(mi_rx_completion_ram_read_data1[143:0])
   ,.mi_rx_completion_ram_read_enable1(mi_rx_completion_ram_read_enable1[1:0])
   ,.mi_rx_completion_ram_err_cor(mi_rx_completion_ram_err_cor[11:0])
   ,.mi_rx_completion_ram_err_uncor(mi_rx_completion_ram_err_uncor[11:0])
   ,.pipe_rx00_char_is_k(pipe_rx00_char_is_k[1:0])
   ,.pipe_rx01_char_is_k(pipe_rx01_char_is_k[1:0])
   ,.pipe_rx02_char_is_k(pipe_rx02_char_is_k[1:0])
   ,.pipe_rx03_char_is_k(pipe_rx03_char_is_k[1:0])
   ,.pipe_rx04_char_is_k(pipe_rx04_char_is_k[1:0])
   ,.pipe_rx05_char_is_k(pipe_rx05_char_is_k[1:0])
   ,.pipe_rx06_char_is_k(pipe_rx06_char_is_k[1:0])
   ,.pipe_rx07_char_is_k(pipe_rx07_char_is_k[1:0])
   ,.pipe_rx08_char_is_k(pipe_rx08_char_is_k[1:0])
   ,.pipe_rx09_char_is_k(pipe_rx09_char_is_k[1:0])
   ,.pipe_rx10_char_is_k(pipe_rx10_char_is_k[1:0])
   ,.pipe_rx11_char_is_k(pipe_rx11_char_is_k[1:0])
   ,.pipe_rx12_char_is_k(pipe_rx12_char_is_k[1:0])
   ,.pipe_rx13_char_is_k(pipe_rx13_char_is_k[1:0])
   ,.pipe_rx14_char_is_k(pipe_rx14_char_is_k[1:0])
   ,.pipe_rx15_char_is_k(pipe_rx15_char_is_k[1:0])
   ,.pipe_rx00_valid(pipe_rx00_valid)
   ,.pipe_rx01_valid(pipe_rx01_valid)
   ,.pipe_rx02_valid(pipe_rx02_valid)
   ,.pipe_rx03_valid(pipe_rx03_valid)
   ,.pipe_rx04_valid(pipe_rx04_valid)
   ,.pipe_rx05_valid(pipe_rx05_valid)
   ,.pipe_rx06_valid(pipe_rx06_valid)
   ,.pipe_rx07_valid(pipe_rx07_valid)
   ,.pipe_rx08_valid(pipe_rx08_valid)
   ,.pipe_rx09_valid(pipe_rx09_valid)
   ,.pipe_rx10_valid(pipe_rx10_valid)
   ,.pipe_rx11_valid(pipe_rx11_valid)
   ,.pipe_rx12_valid(pipe_rx12_valid)
   ,.pipe_rx13_valid(pipe_rx13_valid)
   ,.pipe_rx14_valid(pipe_rx14_valid)
   ,.pipe_rx15_valid(pipe_rx15_valid)
   ,.pipe_rx00_data(pipe_rx00_data[31:0])
   ,.pipe_rx01_data(pipe_rx01_data[31:0])
   ,.pipe_rx02_data(pipe_rx02_data[31:0])
   ,.pipe_rx03_data(pipe_rx03_data[31:0])
   ,.pipe_rx04_data(pipe_rx04_data[31:0])
   ,.pipe_rx05_data(pipe_rx05_data[31:0])
   ,.pipe_rx06_data(pipe_rx06_data[31:0])
   ,.pipe_rx07_data(pipe_rx07_data[31:0])
   ,.pipe_rx08_data(pipe_rx08_data[31:0])
   ,.pipe_rx09_data(pipe_rx09_data[31:0])
   ,.pipe_rx10_data(pipe_rx10_data[31:0])
   ,.pipe_rx11_data(pipe_rx11_data[31:0])
   ,.pipe_rx12_data(pipe_rx12_data[31:0])
   ,.pipe_rx13_data(pipe_rx13_data[31:0])
   ,.pipe_rx14_data(pipe_rx14_data[31:0])
   ,.pipe_rx15_data(pipe_rx15_data[31:0])
   ,.pipe_rx00_polarity(pipe_rx00_polarity)
   ,.pipe_rx01_polarity(pipe_rx01_polarity)
   ,.pipe_rx02_polarity(pipe_rx02_polarity)
   ,.pipe_rx03_polarity(pipe_rx03_polarity)
   ,.pipe_rx04_polarity(pipe_rx04_polarity)
   ,.pipe_rx05_polarity(pipe_rx05_polarity)
   ,.pipe_rx06_polarity(pipe_rx06_polarity)
   ,.pipe_rx07_polarity(pipe_rx07_polarity)
   ,.pipe_rx08_polarity(pipe_rx08_polarity)
   ,.pipe_rx09_polarity(pipe_rx09_polarity)
   ,.pipe_rx10_polarity(pipe_rx10_polarity)
   ,.pipe_rx11_polarity(pipe_rx11_polarity)
   ,.pipe_rx12_polarity(pipe_rx12_polarity)
   ,.pipe_rx13_polarity(pipe_rx13_polarity)
   ,.pipe_rx14_polarity(pipe_rx14_polarity)
   ,.pipe_rx15_polarity(pipe_rx15_polarity)
   ,.pipe_rx00_status(pipe_rx00_status[2:0])
   ,.pipe_rx01_status(pipe_rx01_status[2:0])
   ,.pipe_rx02_status(pipe_rx02_status[2:0])
   ,.pipe_rx03_status(pipe_rx03_status[2:0])
   ,.pipe_rx04_status(pipe_rx04_status[2:0])
   ,.pipe_rx05_status(pipe_rx05_status[2:0])
   ,.pipe_rx06_status(pipe_rx06_status[2:0])
   ,.pipe_rx07_status(pipe_rx07_status[2:0])
   ,.pipe_rx08_status(pipe_rx08_status[2:0])
   ,.pipe_rx09_status(pipe_rx09_status[2:0])
   ,.pipe_rx10_status(pipe_rx10_status[2:0])
   ,.pipe_rx11_status(pipe_rx11_status[2:0])
   ,.pipe_rx12_status(pipe_rx12_status[2:0])
   ,.pipe_rx13_status(pipe_rx13_status[2:0])
   ,.pipe_rx14_status(pipe_rx14_status[2:0])
   ,.pipe_rx15_status(pipe_rx15_status[2:0])
   ,.pipe_rx00_phy_status(pipe_rx00_phy_status)
   ,.pipe_rx01_phy_status(pipe_rx01_phy_status)
   ,.pipe_rx02_phy_status(pipe_rx02_phy_status)
   ,.pipe_rx03_phy_status(pipe_rx03_phy_status)
   ,.pipe_rx04_phy_status(pipe_rx04_phy_status)
   ,.pipe_rx05_phy_status(pipe_rx05_phy_status)
   ,.pipe_rx06_phy_status(pipe_rx06_phy_status)
   ,.pipe_rx07_phy_status(pipe_rx07_phy_status)
   ,.pipe_rx08_phy_status(pipe_rx08_phy_status)
   ,.pipe_rx09_phy_status(pipe_rx09_phy_status)
   ,.pipe_rx10_phy_status(pipe_rx10_phy_status)
   ,.pipe_rx11_phy_status(pipe_rx11_phy_status)
   ,.pipe_rx12_phy_status(pipe_rx12_phy_status)
   ,.pipe_rx13_phy_status(pipe_rx13_phy_status)
   ,.pipe_rx14_phy_status(pipe_rx14_phy_status)
   ,.pipe_rx15_phy_status(pipe_rx15_phy_status)
   ,.pipe_rx00_elec_idle(pipe_rx00_elec_idle)
   ,.pipe_rx01_elec_idle(pipe_rx01_elec_idle)
   ,.pipe_rx02_elec_idle(pipe_rx02_elec_idle)
   ,.pipe_rx03_elec_idle(pipe_rx03_elec_idle)
   ,.pipe_rx04_elec_idle(pipe_rx04_elec_idle)
   ,.pipe_rx05_elec_idle(pipe_rx05_elec_idle)
   ,.pipe_rx06_elec_idle(pipe_rx06_elec_idle)
   ,.pipe_rx07_elec_idle(pipe_rx07_elec_idle)
   ,.pipe_rx08_elec_idle(pipe_rx08_elec_idle)
   ,.pipe_rx09_elec_idle(pipe_rx09_elec_idle)
   ,.pipe_rx10_elec_idle(pipe_rx10_elec_idle)
   ,.pipe_rx11_elec_idle(pipe_rx11_elec_idle)
   ,.pipe_rx12_elec_idle(pipe_rx12_elec_idle)
   ,.pipe_rx13_elec_idle(pipe_rx13_elec_idle)
   ,.pipe_rx14_elec_idle(pipe_rx14_elec_idle)
   ,.pipe_rx15_elec_idle(pipe_rx15_elec_idle)
   ,.pipe_rx00_data_valid(pipe_rx00_data_valid)
   ,.pipe_rx01_data_valid(pipe_rx01_data_valid)
   ,.pipe_rx02_data_valid(pipe_rx02_data_valid)
   ,.pipe_rx03_data_valid(pipe_rx03_data_valid)
   ,.pipe_rx04_data_valid(pipe_rx04_data_valid)
   ,.pipe_rx05_data_valid(pipe_rx05_data_valid)
   ,.pipe_rx06_data_valid(pipe_rx06_data_valid)
   ,.pipe_rx07_data_valid(pipe_rx07_data_valid)
   ,.pipe_rx08_data_valid(pipe_rx08_data_valid)
   ,.pipe_rx09_data_valid(pipe_rx09_data_valid)
   ,.pipe_rx10_data_valid(pipe_rx10_data_valid)
   ,.pipe_rx11_data_valid(pipe_rx11_data_valid)
   ,.pipe_rx12_data_valid(pipe_rx12_data_valid)
   ,.pipe_rx13_data_valid(pipe_rx13_data_valid)
   ,.pipe_rx14_data_valid(pipe_rx14_data_valid)
   ,.pipe_rx15_data_valid(pipe_rx15_data_valid)
   ,.pipe_rx00_start_block(pipe_rx00_start_block[1:0])
   ,.pipe_rx01_start_block(pipe_rx01_start_block[1:0])
   ,.pipe_rx02_start_block(pipe_rx02_start_block[1:0])
   ,.pipe_rx03_start_block(pipe_rx03_start_block[1:0])
   ,.pipe_rx04_start_block(pipe_rx04_start_block[1:0])
   ,.pipe_rx05_start_block(pipe_rx05_start_block[1:0])
   ,.pipe_rx06_start_block(pipe_rx06_start_block[1:0])
   ,.pipe_rx07_start_block(pipe_rx07_start_block[1:0])
   ,.pipe_rx08_start_block(pipe_rx08_start_block[1:0])
   ,.pipe_rx09_start_block(pipe_rx09_start_block[1:0])
   ,.pipe_rx10_start_block(pipe_rx10_start_block[1:0])
   ,.pipe_rx11_start_block(pipe_rx11_start_block[1:0])
   ,.pipe_rx12_start_block(pipe_rx12_start_block[1:0])
   ,.pipe_rx13_start_block(pipe_rx13_start_block[1:0])
   ,.pipe_rx14_start_block(pipe_rx14_start_block[1:0])
   ,.pipe_rx15_start_block(pipe_rx15_start_block[1:0])
   ,.pipe_rx00_sync_header(pipe_rx00_sync_header[1:0])
   ,.pipe_rx01_sync_header(pipe_rx01_sync_header[1:0])
   ,.pipe_rx02_sync_header(pipe_rx02_sync_header[1:0])
   ,.pipe_rx03_sync_header(pipe_rx03_sync_header[1:0])
   ,.pipe_rx04_sync_header(pipe_rx04_sync_header[1:0])
   ,.pipe_rx05_sync_header(pipe_rx05_sync_header[1:0])
   ,.pipe_rx06_sync_header(pipe_rx06_sync_header[1:0])
   ,.pipe_rx07_sync_header(pipe_rx07_sync_header[1:0])
   ,.pipe_rx08_sync_header(pipe_rx08_sync_header[1:0])
   ,.pipe_rx09_sync_header(pipe_rx09_sync_header[1:0])
   ,.pipe_rx10_sync_header(pipe_rx10_sync_header[1:0])
   ,.pipe_rx11_sync_header(pipe_rx11_sync_header[1:0])
   ,.pipe_rx12_sync_header(pipe_rx12_sync_header[1:0])
   ,.pipe_rx13_sync_header(pipe_rx13_sync_header[1:0])
   ,.pipe_rx14_sync_header(pipe_rx14_sync_header[1:0])
   ,.pipe_rx15_sync_header(pipe_rx15_sync_header[1:0])
   ,.pipe_tx00_compliance(pipe_tx00_compliance)
   ,.pipe_tx01_compliance(pipe_tx01_compliance)
   ,.pipe_tx02_compliance(pipe_tx02_compliance)
   ,.pipe_tx03_compliance(pipe_tx03_compliance)
   ,.pipe_tx04_compliance(pipe_tx04_compliance)
   ,.pipe_tx05_compliance(pipe_tx05_compliance)
   ,.pipe_tx06_compliance(pipe_tx06_compliance)
   ,.pipe_tx07_compliance(pipe_tx07_compliance)
   ,.pipe_tx08_compliance(pipe_tx08_compliance)
   ,.pipe_tx09_compliance(pipe_tx09_compliance)
   ,.pipe_tx10_compliance(pipe_tx10_compliance)
   ,.pipe_tx11_compliance(pipe_tx11_compliance)
   ,.pipe_tx12_compliance(pipe_tx12_compliance)
   ,.pipe_tx13_compliance(pipe_tx13_compliance)
   ,.pipe_tx14_compliance(pipe_tx14_compliance)
   ,.pipe_tx15_compliance(pipe_tx15_compliance)
   ,.pipe_tx00_char_is_k(pipe_tx00_char_is_k[1:0])
   ,.pipe_tx01_char_is_k(pipe_tx01_char_is_k[1:0])
   ,.pipe_tx02_char_is_k(pipe_tx02_char_is_k[1:0])
   ,.pipe_tx03_char_is_k(pipe_tx03_char_is_k[1:0])
   ,.pipe_tx04_char_is_k(pipe_tx04_char_is_k[1:0])
   ,.pipe_tx05_char_is_k(pipe_tx05_char_is_k[1:0])
   ,.pipe_tx06_char_is_k(pipe_tx06_char_is_k[1:0])
   ,.pipe_tx07_char_is_k(pipe_tx07_char_is_k[1:0])
   ,.pipe_tx08_char_is_k(pipe_tx08_char_is_k[1:0])
   ,.pipe_tx09_char_is_k(pipe_tx09_char_is_k[1:0])
   ,.pipe_tx10_char_is_k(pipe_tx10_char_is_k[1:0])
   ,.pipe_tx11_char_is_k(pipe_tx11_char_is_k[1:0])
   ,.pipe_tx12_char_is_k(pipe_tx12_char_is_k[1:0])
   ,.pipe_tx13_char_is_k(pipe_tx13_char_is_k[1:0])
   ,.pipe_tx14_char_is_k(pipe_tx14_char_is_k[1:0])
   ,.pipe_tx15_char_is_k(pipe_tx15_char_is_k[1:0])
   ,.pipe_tx00_data(pipe_tx00_data[31:0])
   ,.pipe_tx01_data(pipe_tx01_data[31:0])
   ,.pipe_tx02_data(pipe_tx02_data[31:0])
   ,.pipe_tx03_data(pipe_tx03_data[31:0])
   ,.pipe_tx04_data(pipe_tx04_data[31:0])
   ,.pipe_tx05_data(pipe_tx05_data[31:0])
   ,.pipe_tx06_data(pipe_tx06_data[31:0])
   ,.pipe_tx07_data(pipe_tx07_data[31:0])
   ,.pipe_tx08_data(pipe_tx08_data[31:0])
   ,.pipe_tx09_data(pipe_tx09_data[31:0])
   ,.pipe_tx10_data(pipe_tx10_data[31:0])
   ,.pipe_tx11_data(pipe_tx11_data[31:0])
   ,.pipe_tx12_data(pipe_tx12_data[31:0])
   ,.pipe_tx13_data(pipe_tx13_data[31:0])
   ,.pipe_tx14_data(pipe_tx14_data[31:0])
   ,.pipe_tx15_data(pipe_tx15_data[31:0])
   ,.pipe_tx00_elec_idle(pipe_tx00_elec_idle)
   ,.pipe_tx01_elec_idle(pipe_tx01_elec_idle)
   ,.pipe_tx02_elec_idle(pipe_tx02_elec_idle)
   ,.pipe_tx03_elec_idle(pipe_tx03_elec_idle)
   ,.pipe_tx04_elec_idle(pipe_tx04_elec_idle)
   ,.pipe_tx05_elec_idle(pipe_tx05_elec_idle)
   ,.pipe_tx06_elec_idle(pipe_tx06_elec_idle)
   ,.pipe_tx07_elec_idle(pipe_tx07_elec_idle)
   ,.pipe_tx08_elec_idle(pipe_tx08_elec_idle)
   ,.pipe_tx09_elec_idle(pipe_tx09_elec_idle)
   ,.pipe_tx10_elec_idle(pipe_tx10_elec_idle)
   ,.pipe_tx11_elec_idle(pipe_tx11_elec_idle)
   ,.pipe_tx12_elec_idle(pipe_tx12_elec_idle)
   ,.pipe_tx13_elec_idle(pipe_tx13_elec_idle)
   ,.pipe_tx14_elec_idle(pipe_tx14_elec_idle)
   ,.pipe_tx15_elec_idle(pipe_tx15_elec_idle)
   ,.pipe_tx00_powerdown(pipe_tx00_powerdown[1:0])
   ,.pipe_tx01_powerdown(pipe_tx01_powerdown[1:0])
   ,.pipe_tx02_powerdown(pipe_tx02_powerdown[1:0])
   ,.pipe_tx03_powerdown(pipe_tx03_powerdown[1:0])
   ,.pipe_tx04_powerdown(pipe_tx04_powerdown[1:0])
   ,.pipe_tx05_powerdown(pipe_tx05_powerdown[1:0])
   ,.pipe_tx06_powerdown(pipe_tx06_powerdown[1:0])
   ,.pipe_tx07_powerdown(pipe_tx07_powerdown[1:0])
   ,.pipe_tx08_powerdown(pipe_tx08_powerdown[1:0])
   ,.pipe_tx09_powerdown(pipe_tx09_powerdown[1:0])
   ,.pipe_tx10_powerdown(pipe_tx10_powerdown[1:0])
   ,.pipe_tx11_powerdown(pipe_tx11_powerdown[1:0])
   ,.pipe_tx12_powerdown(pipe_tx12_powerdown[1:0])
   ,.pipe_tx13_powerdown(pipe_tx13_powerdown[1:0])
   ,.pipe_tx14_powerdown(pipe_tx14_powerdown[1:0])
   ,.pipe_tx15_powerdown(pipe_tx15_powerdown[1:0])
   ,.pipe_tx00_data_valid(pipe_tx00_data_valid)
   ,.pipe_tx01_data_valid(pipe_tx01_data_valid)
   ,.pipe_tx02_data_valid(pipe_tx02_data_valid)
   ,.pipe_tx03_data_valid(pipe_tx03_data_valid)
   ,.pipe_tx04_data_valid(pipe_tx04_data_valid)
   ,.pipe_tx05_data_valid(pipe_tx05_data_valid)
   ,.pipe_tx06_data_valid(pipe_tx06_data_valid)
   ,.pipe_tx07_data_valid(pipe_tx07_data_valid)
   ,.pipe_tx08_data_valid(pipe_tx08_data_valid)
   ,.pipe_tx09_data_valid(pipe_tx09_data_valid)
   ,.pipe_tx10_data_valid(pipe_tx10_data_valid)
   ,.pipe_tx11_data_valid(pipe_tx11_data_valid)
   ,.pipe_tx12_data_valid(pipe_tx12_data_valid)
   ,.pipe_tx13_data_valid(pipe_tx13_data_valid)
   ,.pipe_tx14_data_valid(pipe_tx14_data_valid)
   ,.pipe_tx15_data_valid(pipe_tx15_data_valid)
   ,.pipe_tx00_start_block(pipe_tx00_start_block)
   ,.pipe_tx01_start_block(pipe_tx01_start_block)
   ,.pipe_tx02_start_block(pipe_tx02_start_block)
   ,.pipe_tx03_start_block(pipe_tx03_start_block)
   ,.pipe_tx04_start_block(pipe_tx04_start_block)
   ,.pipe_tx05_start_block(pipe_tx05_start_block)
   ,.pipe_tx06_start_block(pipe_tx06_start_block)
   ,.pipe_tx07_start_block(pipe_tx07_start_block)
   ,.pipe_tx08_start_block(pipe_tx08_start_block)
   ,.pipe_tx09_start_block(pipe_tx09_start_block)
   ,.pipe_tx10_start_block(pipe_tx10_start_block)
   ,.pipe_tx11_start_block(pipe_tx11_start_block)
   ,.pipe_tx12_start_block(pipe_tx12_start_block)
   ,.pipe_tx13_start_block(pipe_tx13_start_block)
   ,.pipe_tx14_start_block(pipe_tx14_start_block)
   ,.pipe_tx15_start_block(pipe_tx15_start_block)
   ,.pipe_tx00_sync_header(pipe_tx00_sync_header[1:0])
   ,.pipe_tx01_sync_header(pipe_tx01_sync_header[1:0])
   ,.pipe_tx02_sync_header(pipe_tx02_sync_header[1:0])
   ,.pipe_tx03_sync_header(pipe_tx03_sync_header[1:0])
   ,.pipe_tx04_sync_header(pipe_tx04_sync_header[1:0])
   ,.pipe_tx05_sync_header(pipe_tx05_sync_header[1:0])
   ,.pipe_tx06_sync_header(pipe_tx06_sync_header[1:0])
   ,.pipe_tx07_sync_header(pipe_tx07_sync_header[1:0])
   ,.pipe_tx08_sync_header(pipe_tx08_sync_header[1:0])
   ,.pipe_tx09_sync_header(pipe_tx09_sync_header[1:0])
   ,.pipe_tx10_sync_header(pipe_tx10_sync_header[1:0])
   ,.pipe_tx11_sync_header(pipe_tx11_sync_header[1:0])
   ,.pipe_tx12_sync_header(pipe_tx12_sync_header[1:0])
   ,.pipe_tx13_sync_header(pipe_tx13_sync_header[1:0])
   ,.pipe_tx14_sync_header(pipe_tx14_sync_header[1:0])
   ,.pipe_tx15_sync_header(pipe_tx15_sync_header[1:0])
   ,.pipe_rx00_eq_control(pipe_rx00_eq_control[1:0])
   ,.pipe_rx01_eq_control(pipe_rx01_eq_control[1:0])
   ,.pipe_rx02_eq_control(pipe_rx02_eq_control[1:0])
   ,.pipe_rx03_eq_control(pipe_rx03_eq_control[1:0])
   ,.pipe_rx04_eq_control(pipe_rx04_eq_control[1:0])
   ,.pipe_rx05_eq_control(pipe_rx05_eq_control[1:0])
   ,.pipe_rx06_eq_control(pipe_rx06_eq_control[1:0])
   ,.pipe_rx07_eq_control(pipe_rx07_eq_control[1:0])
   ,.pipe_rx08_eq_control(pipe_rx08_eq_control[1:0])
   ,.pipe_rx09_eq_control(pipe_rx09_eq_control[1:0])
   ,.pipe_rx10_eq_control(pipe_rx10_eq_control[1:0])
   ,.pipe_rx11_eq_control(pipe_rx11_eq_control[1:0])
   ,.pipe_rx12_eq_control(pipe_rx12_eq_control[1:0])
   ,.pipe_rx13_eq_control(pipe_rx13_eq_control[1:0])
   ,.pipe_rx14_eq_control(pipe_rx14_eq_control[1:0])
   ,.pipe_rx15_eq_control(pipe_rx15_eq_control[1:0])
   ,.pipe_rx00_eq_lp_lf_fs_sel(pipe_rx00_eq_lp_lf_fs_sel)
   ,.pipe_rx01_eq_lp_lf_fs_sel(pipe_rx01_eq_lp_lf_fs_sel)
   ,.pipe_rx02_eq_lp_lf_fs_sel(pipe_rx02_eq_lp_lf_fs_sel)
   ,.pipe_rx03_eq_lp_lf_fs_sel(pipe_rx03_eq_lp_lf_fs_sel)
   ,.pipe_rx04_eq_lp_lf_fs_sel(pipe_rx04_eq_lp_lf_fs_sel)
   ,.pipe_rx05_eq_lp_lf_fs_sel(pipe_rx05_eq_lp_lf_fs_sel)
   ,.pipe_rx06_eq_lp_lf_fs_sel(pipe_rx06_eq_lp_lf_fs_sel)
   ,.pipe_rx07_eq_lp_lf_fs_sel(pipe_rx07_eq_lp_lf_fs_sel)
   ,.pipe_rx08_eq_lp_lf_fs_sel(pipe_rx08_eq_lp_lf_fs_sel)
   ,.pipe_rx09_eq_lp_lf_fs_sel(pipe_rx09_eq_lp_lf_fs_sel)
   ,.pipe_rx10_eq_lp_lf_fs_sel(pipe_rx10_eq_lp_lf_fs_sel)
   ,.pipe_rx11_eq_lp_lf_fs_sel(pipe_rx11_eq_lp_lf_fs_sel)
   ,.pipe_rx12_eq_lp_lf_fs_sel(pipe_rx12_eq_lp_lf_fs_sel)
   ,.pipe_rx13_eq_lp_lf_fs_sel(pipe_rx13_eq_lp_lf_fs_sel)
   ,.pipe_rx14_eq_lp_lf_fs_sel(pipe_rx14_eq_lp_lf_fs_sel)
   ,.pipe_rx15_eq_lp_lf_fs_sel(pipe_rx15_eq_lp_lf_fs_sel)
   ,.pipe_rx00_eq_lp_new_tx_coeff_or_preset(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx01_eq_lp_new_tx_coeff_or_preset(pipe_rx01_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx02_eq_lp_new_tx_coeff_or_preset(pipe_rx02_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx03_eq_lp_new_tx_coeff_or_preset(pipe_rx03_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx04_eq_lp_new_tx_coeff_or_preset(pipe_rx04_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx05_eq_lp_new_tx_coeff_or_preset(pipe_rx05_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx06_eq_lp_new_tx_coeff_or_preset(pipe_rx06_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx07_eq_lp_new_tx_coeff_or_preset(pipe_rx07_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx08_eq_lp_new_tx_coeff_or_preset(pipe_rx08_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx09_eq_lp_new_tx_coeff_or_preset(pipe_rx09_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx10_eq_lp_new_tx_coeff_or_preset(pipe_rx10_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx11_eq_lp_new_tx_coeff_or_preset(pipe_rx11_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx12_eq_lp_new_tx_coeff_or_preset(pipe_rx12_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx13_eq_lp_new_tx_coeff_or_preset(pipe_rx13_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx14_eq_lp_new_tx_coeff_or_preset(pipe_rx14_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx15_eq_lp_new_tx_coeff_or_preset(pipe_rx15_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.pipe_rx00_eq_lp_adapt_done(pipe_rx00_eq_lp_adapt_done)
   ,.pipe_rx01_eq_lp_adapt_done(pipe_rx01_eq_lp_adapt_done)
   ,.pipe_rx02_eq_lp_adapt_done(pipe_rx02_eq_lp_adapt_done)
   ,.pipe_rx03_eq_lp_adapt_done(pipe_rx03_eq_lp_adapt_done)
   ,.pipe_rx04_eq_lp_adapt_done(pipe_rx04_eq_lp_adapt_done)
   ,.pipe_rx05_eq_lp_adapt_done(pipe_rx05_eq_lp_adapt_done)
   ,.pipe_rx06_eq_lp_adapt_done(pipe_rx06_eq_lp_adapt_done)
   ,.pipe_rx07_eq_lp_adapt_done(pipe_rx07_eq_lp_adapt_done)
   ,.pipe_rx08_eq_lp_adapt_done(pipe_rx08_eq_lp_adapt_done)
   ,.pipe_rx09_eq_lp_adapt_done(pipe_rx09_eq_lp_adapt_done)
   ,.pipe_rx10_eq_lp_adapt_done(pipe_rx10_eq_lp_adapt_done)
   ,.pipe_rx11_eq_lp_adapt_done(pipe_rx11_eq_lp_adapt_done)
   ,.pipe_rx12_eq_lp_adapt_done(pipe_rx12_eq_lp_adapt_done)
   ,.pipe_rx13_eq_lp_adapt_done(pipe_rx13_eq_lp_adapt_done)
   ,.pipe_rx14_eq_lp_adapt_done(pipe_rx14_eq_lp_adapt_done)
   ,.pipe_rx15_eq_lp_adapt_done(pipe_rx15_eq_lp_adapt_done)
   ,.pipe_rx00_eq_done(pipe_rx00_eq_done)
   ,.pipe_rx01_eq_done(pipe_rx01_eq_done)
   ,.pipe_rx02_eq_done(pipe_rx02_eq_done)
   ,.pipe_rx03_eq_done(pipe_rx03_eq_done)
   ,.pipe_rx04_eq_done(pipe_rx04_eq_done)
   ,.pipe_rx05_eq_done(pipe_rx05_eq_done)
   ,.pipe_rx06_eq_done(pipe_rx06_eq_done)
   ,.pipe_rx07_eq_done(pipe_rx07_eq_done)
   ,.pipe_rx08_eq_done(pipe_rx08_eq_done)
   ,.pipe_rx09_eq_done(pipe_rx09_eq_done)
   ,.pipe_rx10_eq_done(pipe_rx10_eq_done)
   ,.pipe_rx11_eq_done(pipe_rx11_eq_done)
   ,.pipe_rx12_eq_done(pipe_rx12_eq_done)
   ,.pipe_rx13_eq_done(pipe_rx13_eq_done)
   ,.pipe_rx14_eq_done(pipe_rx14_eq_done)
   ,.pipe_rx15_eq_done(pipe_rx15_eq_done)
   ,.pipe_tx00_eq_control(pipe_tx00_eq_control[1:0])
   ,.pipe_tx01_eq_control(pipe_tx01_eq_control[1:0])
   ,.pipe_tx02_eq_control(pipe_tx02_eq_control[1:0])
   ,.pipe_tx03_eq_control(pipe_tx03_eq_control[1:0])
   ,.pipe_tx04_eq_control(pipe_tx04_eq_control[1:0])
   ,.pipe_tx05_eq_control(pipe_tx05_eq_control[1:0])
   ,.pipe_tx06_eq_control(pipe_tx06_eq_control[1:0])
   ,.pipe_tx07_eq_control(pipe_tx07_eq_control[1:0])
   ,.pipe_tx08_eq_control(pipe_tx08_eq_control[1:0])
   ,.pipe_tx09_eq_control(pipe_tx09_eq_control[1:0])
   ,.pipe_tx10_eq_control(pipe_tx10_eq_control[1:0])
   ,.pipe_tx11_eq_control(pipe_tx11_eq_control[1:0])
   ,.pipe_tx12_eq_control(pipe_tx12_eq_control[1:0])
   ,.pipe_tx13_eq_control(pipe_tx13_eq_control[1:0])
   ,.pipe_tx14_eq_control(pipe_tx14_eq_control[1:0])
   ,.pipe_tx15_eq_control(pipe_tx15_eq_control[1:0])
   ,.pipe_tx00_eq_deemph(pipe_tx00_eq_deemph[5:0])
   ,.pipe_tx01_eq_deemph(pipe_tx01_eq_deemph[5:0])
   ,.pipe_tx02_eq_deemph(pipe_tx02_eq_deemph[5:0])
   ,.pipe_tx03_eq_deemph(pipe_tx03_eq_deemph[5:0])
   ,.pipe_tx04_eq_deemph(pipe_tx04_eq_deemph[5:0])
   ,.pipe_tx05_eq_deemph(pipe_tx05_eq_deemph[5:0])
   ,.pipe_tx06_eq_deemph(pipe_tx06_eq_deemph[5:0])
   ,.pipe_tx07_eq_deemph(pipe_tx07_eq_deemph[5:0])
   ,.pipe_tx08_eq_deemph(pipe_tx08_eq_deemph[5:0])
   ,.pipe_tx09_eq_deemph(pipe_tx09_eq_deemph[5:0])
   ,.pipe_tx10_eq_deemph(pipe_tx10_eq_deemph[5:0])
   ,.pipe_tx11_eq_deemph(pipe_tx11_eq_deemph[5:0])
   ,.pipe_tx12_eq_deemph(pipe_tx12_eq_deemph[5:0])
   ,.pipe_tx13_eq_deemph(pipe_tx13_eq_deemph[5:0])
   ,.pipe_tx14_eq_deemph(pipe_tx14_eq_deemph[5:0])
   ,.pipe_tx15_eq_deemph(pipe_tx15_eq_deemph[5:0])
   ,.pipe_tx00_eq_coeff(pipe_tx00_eq_coeff[17:0])
   ,.pipe_tx01_eq_coeff(pipe_tx01_eq_coeff[17:0])
   ,.pipe_tx02_eq_coeff(pipe_tx02_eq_coeff[17:0])
   ,.pipe_tx03_eq_coeff(pipe_tx03_eq_coeff[17:0])
   ,.pipe_tx04_eq_coeff(pipe_tx04_eq_coeff[17:0])
   ,.pipe_tx05_eq_coeff(pipe_tx05_eq_coeff[17:0])
   ,.pipe_tx06_eq_coeff(pipe_tx06_eq_coeff[17:0])
   ,.pipe_tx07_eq_coeff(pipe_tx07_eq_coeff[17:0])
   ,.pipe_tx08_eq_coeff(pipe_tx08_eq_coeff[17:0])
   ,.pipe_tx09_eq_coeff(pipe_tx09_eq_coeff[17:0])
   ,.pipe_tx10_eq_coeff(pipe_tx10_eq_coeff[17:0])
   ,.pipe_tx11_eq_coeff(pipe_tx11_eq_coeff[17:0])
   ,.pipe_tx12_eq_coeff(pipe_tx12_eq_coeff[17:0])
   ,.pipe_tx13_eq_coeff(pipe_tx13_eq_coeff[17:0])
   ,.pipe_tx14_eq_coeff(pipe_tx14_eq_coeff[17:0])
   ,.pipe_tx15_eq_coeff(pipe_tx15_eq_coeff[17:0])
   ,.pipe_tx00_eq_done(pipe_tx00_eq_done)
   ,.pipe_tx01_eq_done(pipe_tx01_eq_done)
   ,.pipe_tx02_eq_done(pipe_tx02_eq_done)
   ,.pipe_tx03_eq_done(pipe_tx03_eq_done)
   ,.pipe_tx04_eq_done(pipe_tx04_eq_done)
   ,.pipe_tx05_eq_done(pipe_tx05_eq_done)
   ,.pipe_tx06_eq_done(pipe_tx06_eq_done)
   ,.pipe_tx07_eq_done(pipe_tx07_eq_done)
   ,.pipe_tx08_eq_done(pipe_tx08_eq_done)
   ,.pipe_tx09_eq_done(pipe_tx09_eq_done)
   ,.pipe_tx10_eq_done(pipe_tx10_eq_done)
   ,.pipe_tx11_eq_done(pipe_tx11_eq_done)
   ,.pipe_tx12_eq_done(pipe_tx12_eq_done)
   ,.pipe_tx13_eq_done(pipe_tx13_eq_done)
   ,.pipe_tx14_eq_done(pipe_tx14_eq_done)
   ,.pipe_tx15_eq_done(pipe_tx15_eq_done)
   ,.pipe_rx_eq_lp_tx_preset(pipe_rx_eq_lp_tx_preset[3:0])
   ,.pipe_rx_eq_lp_lf_fs(pipe_rx_eq_lp_lf_fs[5:0])
   ,.pipe_tx_rcvr_det(pipe_tx_rcvr_det)
   ,.pipe_tx_rate(pipe_tx_rate[1:0])
   ,.pipe_tx_deemph(pipe_tx_deemph)
   ,.pipe_tx_margin(pipe_tx_margin[2:0])
   ,.pipe_tx_swing(pipe_tx_swing)
   ,.pipe_tx_reset(pipe_tx_reset)
   ,.pipe_eq_fs(pipe_eq_fs[5:0])
   ,.pipe_eq_lf(pipe_eq_lf[5:0])
   ,.pl_gen2_upstream_prefer_deemph(pl_gen2_upstream_prefer_deemph)
   ,.pl_eq_in_progress(pl_eq_in_progress)
   ,.pl_eq_phase(pl_eq_phase[1:0])
   ,.pl_eq_reset_eieos_count(pl_eq_reset_eieos_count)
   ,.pl_gen34_redo_equalization(pl_gen34_redo_equalization)
   ,.pl_gen34_redo_eq_speed(pl_gen34_redo_eq_speed)
   ,.pl_gen34_eq_mismatch(pl_gen34_eq_mismatch)
   ,.m_axis_cq_tdata(m_axis_cq_tdata_int[255:0])
   ,.s_axis_cc_tdata(s_axis_cc_tdata_int[255:0])
   ,.s_axis_rq_tdata(s_axis_rq_tdata_int[255:0])
   ,.m_axis_rc_tdata(m_axis_rc_tdata_int[255:0])
   ,.m_axis_cq_tuser(m_axis_cq_tuser_int[87:0])
   ,.s_axis_cc_tuser(s_axis_cc_tuser_int[32:0])
   ,.m_axis_cq_tlast(m_axis_cq_tlast_int)
   ,.s_axis_rq_tlast(s_axis_rq_tlast_int)
   ,.m_axis_rc_tlast(m_axis_rc_tlast_int)
   ,.s_axis_cc_tlast(s_axis_cc_tlast_int)
   ,.pcie_cq_np_req(pcie_cq_np_req[1:0])
   ,.pcie_cq_np_req_count(pcie_cq_np_req_count_int[5:0])
   ,.s_axis_rq_tuser(s_axis_rq_tuser_int[61:0])
   ,.m_axis_rc_tuser(m_axis_rc_tuser_int[74:0])
   ,.m_axis_cq_tkeep(m_axis_cq_tkeep_int[7:0])
   ,.s_axis_cc_tkeep(s_axis_cc_tkeep_int[7:0])
   ,.s_axis_rq_tkeep(s_axis_rq_tkeep_int[7:0])
   ,.m_axis_rc_tkeep(m_axis_rc_tkeep_int[7:0])
   ,.m_axis_cq_tvalid(m_axis_cq_tvalid_int)
   ,.s_axis_cc_tvalid(s_axis_cc_tvalid_int)
   ,.s_axis_rq_tvalid(s_axis_rq_tvalid_int)
   ,.m_axis_rc_tvalid(m_axis_rc_tvalid_int)
   ,.m_axis_cq_tready(m_axis_cq_tready_int[21:0])
   ,.s_axis_cc_tready(s_axis_cc_tready_int[3:0])
   ,.s_axis_rq_tready(s_axis_rq_tready_int[3:0])
   ,.m_axis_rc_tready(m_axis_rc_tready_int[21:0])
   ,.pcie_rq_seq_num0(pcie_rq_seq_num0_cc[5:0])
   ,.pcie_rq_seq_num_vld0(pcie_rq_seq_num_vld0_cc)
   ,.pcie_rq_seq_num1(pcie_rq_seq_num1[5:0])
   ,.pcie_rq_seq_num_vld1(pcie_rq_seq_num_vld1)
   ,.pcie_rq_tag0(pcie_rq_tag0[7:0])
   ,.pcie_rq_tag_vld0(pcie_rq_tag_vld0)
   ,.pcie_rq_tag1(pcie_rq_tag1[7:0])
   ,.pcie_rq_tag_vld1(pcie_rq_tag_vld1)
   ,.pcie_tfc_nph_av(pcie_tfc_nph_av[3:0])
   ,.pcie_tfc_npd_av(pcie_tfc_npd_av[3:0])
   ,.pcie_rq_tag_av(pcie_rq_tag_av[3:0])
   ,.pcie_posted_req_delivered(pcie_posted_req_delivered)
   ,.pcie_cq_pipeline_empty(pcie_cq_pipeline_empty)
   ,.pcie_cq_np_user_credit_rcvd(pcie_cq_np_user_credit_rcvd)
   ,.pcie_compl_delivered(pcie_compl_delivered[1:0])
   ,.pcie_compl_delivered_tag0(pcie_compl_delivered_tag0[7:0])
   ,.pcie_compl_delivered_tag1(pcie_compl_delivered_tag1[7:0])
   ,.axi_user_out(axi_user_out[7:0])
   ,.axi_user_in(axi_user_in[7:0])
   ,.cfg_mgmt_addr(cfg_mgmt_addr[9:0])
   ,.cfg_mgmt_function_number(cfg_mgmt_function_number[7:0])
   ,.cfg_mgmt_write(cfg_mgmt_write)
   ,.cfg_mgmt_write_data(cfg_mgmt_write_data[31:0])
   ,.cfg_mgmt_byte_enable(cfg_mgmt_byte_enable[3:0])
   ,.cfg_mgmt_read(cfg_mgmt_read)
   ,.cfg_mgmt_read_data(cfg_mgmt_read_data[31:0])
   ,.cfg_mgmt_read_write_done(cfg_mgmt_read_write_done)
   ,.cfg_mgmt_debug_access(cfg_mgmt_debug_access)
   ,.cfg_phy_link_down(cfg_phy_link_down_wire)
   ,.cfg_phy_link_status(cfg_phy_link_status[1:0])
   ,.cfg_negotiated_width(cfg_negotiated_width[2:0])
   ,.cfg_current_speed(cfg_current_speed[1:0])
   ,.cfg_max_payload(cfg_max_payload[1:0])
   ,.cfg_max_read_req(cfg_max_read_req[2:0])
   ,.cfg_function_status(cfg_function_status[15:0])
   ,.cfg_function_power_state(cfg_function_power_state[11:0])
   ,.cfg_link_power_state(cfg_link_power_state[1:0])
   ,.cfg_err_cor_out(cfg_err_cor_out)
   ,.cfg_err_nonfatal_out(cfg_err_nonfatal_out)
   ,.cfg_err_fatal_out(cfg_err_fatal_out)
   ,.cfg_local_error_valid(cfg_local_error_valid)
   ,.cfg_local_error_out(cfg_local_error_out[4:0])
   ,.cfg_ltr_enable(cfg_ltr_enable)
   ,.cfg_ltssm_state(cfg_ltssm_state[5:0])
   ,.cfg_rx_pm_state(cfg_rx_pm_state[1:0])
   ,.cfg_tx_pm_state(cfg_tx_pm_state[1:0])
   ,.cfg_rcb_status(cfg_rcb_status[3:0])
   ,.cfg_obff_enable(cfg_obff_enable[1:0])
   ,.cfg_pl_status_change(cfg_pl_status_change)
   ,.cfg_tph_requester_enable(cfg_tph_requester_enable[3:0])
   ,.cfg_tph_st_mode(cfg_tph_st_mode[11:0])
   ,.cfg_msg_received(cfg_msg_received)
   ,.cfg_msg_received_data(cfg_msg_received_data[7:0])
   ,.cfg_msg_received_type(cfg_msg_received_type[4:0])
   ,.cfg_msg_transmit(cfg_msg_transmit)
   ,.cfg_msg_transmit_type(cfg_msg_transmit_type[2:0])
   ,.cfg_msg_transmit_data(cfg_msg_transmit_data[31:0])
   ,.cfg_msg_transmit_done(cfg_msg_transmit_done)
   ,.cfg_fc_ph(cfg_fc_ph[7:0])
   ,.cfg_fc_pd(cfg_fc_pd[11:0])
   ,.cfg_fc_nph(cfg_fc_nph[7:0])
   ,.cfg_fc_npd(cfg_fc_npd[11:0])
   ,.cfg_fc_cplh(cfg_fc_cplh[7:0])
   ,.cfg_fc_cpld(cfg_fc_cpld[11:0])
   ,.cfg_fc_sel(cfg_fc_sel[2:0])
   ,.cfg_hot_reset_in(cfg_hot_reset_in)
   ,.cfg_hot_reset_out(cfg_hot_reset_out)
   ,.cfg_config_space_enable(cfg_config_space_enable)
   ,.cfg_dsn(cfg_dsn[63:0])
   ,.cfg_dev_id_pf0(cfg_dev_id_pf0[15:0])
   ,.cfg_dev_id_pf1(cfg_dev_id_pf1[15:0])
   ,.cfg_dev_id_pf2(cfg_dev_id_pf2[15:0])
   ,.cfg_dev_id_pf3(cfg_dev_id_pf3[15:0])
   ,.cfg_vend_id(cfg_vend_id[15:0])
   ,.cfg_rev_id_pf0(cfg_rev_id_pf0[7:0])
   ,.cfg_rev_id_pf1(cfg_rev_id_pf1[7:0])
   ,.cfg_rev_id_pf2(cfg_rev_id_pf2[7:0])
   ,.cfg_rev_id_pf3(cfg_rev_id_pf3[7:0])
   ,.cfg_subsys_id_pf0(cfg_subsys_id_pf0[15:0])
   ,.cfg_subsys_id_pf1(cfg_subsys_id_pf1[15:0])
   ,.cfg_subsys_id_pf2(cfg_subsys_id_pf2[15:0])
   ,.cfg_subsys_id_pf3(cfg_subsys_id_pf3[15:0])
   ,.cfg_subsys_vend_id(cfg_subsys_vend_id[15:0])
   ,.cfg_ds_port_number(cfg_ds_port_number[7:0])
   ,.cfg_ds_bus_number(cfg_ds_bus_number[7:0])
   ,.cfg_ds_device_number(cfg_ds_device_number[4:0])
   ,.cfg_ds_function_number(cfg_ds_function_number[2:0])
   ,.cfg_bus_number(cfg_bus_number[7:0])
   ,.cfg_power_state_change_ack(cfg_power_state_change_ack)
   ,.cfg_power_state_change_interrupt(cfg_power_state_change_interrupt)
   ,.cfg_err_cor_in(cfg_err_cor_in)
   ,.cfg_err_uncor_in(cfg_err_uncor_in)
   ,.cfg_flr_done(cfg_flr_done[3:0])
   ,.cfg_vf_flr_func_num(cfg_vf_flr_func_num[7:0])
   ,.cfg_vf_flr_done(cfg_vf_flr_done)
   ,.cfg_flr_in_process(cfg_flr_in_process[3:0])
   ,.cfg_req_pm_transition_l23_ready(cfg_req_pm_transition_l23_ready)
   ,.cfg_link_training_enable(cfg_link_training_enable)
   ,.cfg_interrupt_int(cfg_interrupt_int[3:0])
   ,.cfg_interrupt_sent(cfg_interrupt_sent)
   ,.cfg_interrupt_pending(cfg_interrupt_pending[3:0])
   ,.cfg_interrupt_msi_enable(cfg_interrupt_msi_enable[3:0])
   ,.cfg_interrupt_msi_int(cfg_interrupt_msi_int[31:0])
   ,.cfg_interrupt_msi_sent(cfg_interrupt_msi_sent)
   ,.cfg_interrupt_msi_fail(cfg_interrupt_msi_fail)
   ,.cfg_interrupt_msi_mmenable(cfg_interrupt_msi_mmenable[11:0])
   ,.cfg_interrupt_msi_pending_status(cfg_interrupt_msi_pending_status[31:0])
   ,.cfg_interrupt_msi_pending_status_function_num(cfg_interrupt_msi_pending_status_function_num[1:0])
   ,.cfg_interrupt_msi_pending_status_data_enable(cfg_interrupt_msi_pending_status_data_enable)
   ,.cfg_interrupt_msi_mask_update(cfg_interrupt_msi_mask_update)
   ,.cfg_interrupt_msi_select(cfg_interrupt_msi_select[1:0])
   ,.cfg_interrupt_msi_data(cfg_interrupt_msi_data[31:0])
   ,.cfg_interrupt_msix_enable(cfg_interrupt_msix_enable[3:0])
   ,.cfg_interrupt_msix_mask(cfg_interrupt_msix_mask[3:0])
   ,.cfg_interrupt_msix_address(cfg_interrupt_msix_address[63:0])
   ,.cfg_interrupt_msix_data(cfg_interrupt_msix_data[31:0])
   ,.cfg_interrupt_msix_int(cfg_interrupt_msix_int)
   ,.cfg_interrupt_msix_vec_pending(cfg_interrupt_msix_vec_pending[1:0])
   ,.cfg_interrupt_msix_vec_pending_status(cfg_interrupt_msix_vec_pending_status)
   ,.cfg_interrupt_msi_attr(cfg_interrupt_msi_attr[2:0])
   ,.cfg_interrupt_msi_tph_present(cfg_interrupt_msi_tph_present)
   ,.cfg_interrupt_msi_tph_type(cfg_interrupt_msi_tph_type[1:0])
   ,.cfg_interrupt_msi_tph_st_tag(cfg_interrupt_msi_tph_st_tag[7:0])
   ,.cfg_interrupt_msi_function_number(cfg_interrupt_msi_function_number[7:0])
   ,.cfg_ext_read_received(cfg_ext_read_received)
   ,.cfg_ext_write_received(cfg_ext_write_received)
   ,.cfg_ext_register_number(cfg_ext_register_number[9:0])
   ,.cfg_ext_function_number(cfg_ext_function_number[7:0])
   ,.cfg_ext_write_data(cfg_ext_write_data[31:0])
   ,.cfg_ext_write_byte_enable(cfg_ext_write_byte_enable[3:0])
   ,.cfg_ext_read_data(cfg_ext_read_data[31:0])
   ,.cfg_ext_read_data_valid(cfg_ext_read_data_valid)
   ,.cfg_tph_ram_address(cfg_tph_ram_address[11:0])
   ,.cfg_tph_ram_write_data(cfg_tph_ram_write_data[35:0])
   ,.cfg_tph_ram_write_byte_enable(cfg_tph_ram_write_byte_enable[3:0])
   ,.cfg_tph_ram_read_data(cfg_tph_ram_read_data[35:0])
   ,.cfg_tph_ram_read_enable(cfg_tph_ram_read_enable)
   ,.cfg_msix_ram_address(cfg_msix_ram_address[12:0])
   ,.cfg_msix_ram_write_data(cfg_msix_ram_write_data[35:0])
   ,.cfg_msix_ram_write_byte_enable(cfg_msix_ram_write_byte_enable[3:0])
   ,.cfg_msix_ram_read_data(cfg_msix_ram_read_data[35:0])
   ,.cfg_msix_ram_read_enable(cfg_msix_ram_read_enable)
   ,.cfg_pm_aspm_l1_entry_reject(cfg_pm_aspm_l1_entry_reject)
   ,.cfg_pm_aspm_tx_l0s_entry_disable(cfg_pm_aspm_tx_l0s_entry_disable)
   ,.conf_req_type(conf_req_type[1:0])
   ,.conf_req_reg_num(conf_req_reg_num[3:0])
   ,.conf_req_data(conf_req_data[31:0])
   ,.conf_req_valid(conf_req_valid)
   ,.conf_req_ready(conf_req_ready)
   ,.conf_resp_rdata(conf_resp_rdata[31:0])
   ,.conf_resp_valid(conf_resp_valid)
   ,.conf_mcap_design_switch(conf_mcap_design_switch)
   ,.conf_mcap_eos(conf_mcap_eos)
   ,.conf_mcap_in_use_by_pcie(conf_mcap_in_use_by_pcie)
   ,.conf_mcap_request_by_conf(conf_mcap_request_by_conf)
   ,.dbg_data0_out( )
   ,.dbg_ctrl0_out( )
   ,.dbg_sel0(6'd0)
   ,.dbg_data1_out( )
   ,.dbg_ctrl1_out( )
   ,.dbg_sel1(6'd0)
   ,.drp_clk(drp_clk)
   ,.drp_en(drp_en)
   ,.drp_we(drp_we)
   ,.drp_addr(drp_addr[9:0])
   ,.drp_di(drp_di[15:0])
   ,.drp_rdy(drp_rdy)
   ,.drp_do(drp_do[15:0])
   ,.scanmode_n(1'b0)
   ,.scanenable_n(1'b0)
   ,.scanin({150{1'b0}})
   ,.scanout( )
   ,.pipe_clk(pipe_clk_to_e4)
   ,.core_clk(core_clk)
   ,.core_clk_mi_replay_ram0(core_clk)
   ,.core_clk_mi_replay_ram1(core_clk)
   ,.core_clk_mi_rx_completion_ram0(core_clk)
   ,.core_clk_mi_rx_completion_ram1(core_clk)
   ,.core_clk_mi_rx_posted_request_ram0(core_clk)
   ,.core_clk_mi_rx_posted_request_ram1(core_clk)
   ,.user_clk(user_clk_to_e4)
   ,.user_clk2(user_clk2_to_e4)
   ,.mcap_clk(mcap_clk)
   ,.mcap_rst_b(mcap_rst_b)
   ,.reset_n(reset_n)
   ,.mgmt_reset_n(mgmt_reset_n)
   ,.mgmt_sticky_reset_n(mgmt_sticky_reset_n)
   ,.pipe_reset_n(pipe_reset_n)
   ,.pcie_perst0_b(pcie_perst0_b)
   ,.pcie_perst1_b(pcie_perst1_b)
   ,.user_clk_en(user_clk_en_to_e4) // note name change
   ,.pipe_clk_en(1'b1)
   ,.pmv_enable_n(1'b0)
   ,.pmv_select(3'b000)
   ,.pmv_divide(2'b00)
   ,.pmv_out( )
   ,.user_spare_in({32{1'b0}})
   ,.user_spare_out( )
  );

  end else begin : pcie_4_0_genblk // IMPL_TARGET == "HARD"

  PCIE40E4 #(

    .CRM_CORE_CLK_FREQ_500(CRM_CORE_CLK_FREQ_500)
   ,.CRM_USER_CLK_FREQ(CRM_USER_CLK_FREQ)
   ,.SIM_DEVICE(SIM_DEVICE)
   ,.AXISTEN_IF_WIDTH(AXISTEN_IF_WIDTH)
   ,.AXISTEN_IF_EXT_512(AXISTEN_IF_EXT_512)
   ,.AXISTEN_IF_EXT_512_CQ_STRADDLE(AXISTEN_IF_EXT_512_CQ_STRADDLE)
   ,.AXISTEN_IF_EXT_512_CC_STRADDLE(AXISTEN_IF_EXT_512_CC_STRADDLE)
   ,.AXISTEN_IF_EXT_512_RQ_STRADDLE(AXISTEN_IF_EXT_512_RQ_STRADDLE)
   ,.AXISTEN_IF_EXT_512_RC_STRADDLE(AXISTEN_IF_EXT_512_RC_STRADDLE)
   ,.AXISTEN_IF_CQ_ALIGNMENT_MODE(AXISTEN_IF_CQ_ALIGNMENT_MODE)
   ,.AXISTEN_IF_CC_ALIGNMENT_MODE(AXISTEN_IF_CC_ALIGNMENT_MODE)
   ,.AXISTEN_IF_RQ_ALIGNMENT_MODE(AXISTEN_IF_RQ_ALIGNMENT_MODE)
   ,.AXISTEN_IF_RC_ALIGNMENT_MODE(AXISTEN_IF_RC_ALIGNMENT_MODE)
   ,.AXISTEN_IF_RC_STRADDLE(AXISTEN_IF_RC_STRADDLE)
   ,.AXISTEN_IF_ENABLE_RX_MSG_INTFC(AXISTEN_IF_ENABLE_RX_MSG_INTFC)
   ,.AXISTEN_IF_ENABLE_MSG_ROUTE(AXISTEN_IF_ENABLE_MSG_ROUTE)
   ,.AXISTEN_IF_RX_PARITY_EN(AXISTEN_IF_RX_PARITY_EN)
   ,.AXISTEN_IF_TX_PARITY_EN(AXISTEN_IF_TX_PARITY_EN)
   ,.AXISTEN_IF_ENABLE_CLIENT_TAG(AXISTEN_IF_ENABLE_CLIENT_TAG)
   ,.AXISTEN_IF_ENABLE_256_TAGS(AXISTEN_IF_ENABLE_256_TAGS)
   ,.AXISTEN_IF_COMPL_TIMEOUT_REG0(AXISTEN_IF_COMPL_TIMEOUT_REG0)
   ,.AXISTEN_IF_COMPL_TIMEOUT_REG1(AXISTEN_IF_COMPL_TIMEOUT_REG1)
   ,.AXISTEN_IF_LEGACY_MODE_ENABLE(AXISTEN_IF_LEGACY_MODE_ENABLE)
   ,.AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK(AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK)
   ,.AXISTEN_IF_MSIX_TO_RAM_PIPELINE(AXISTEN_IF_MSIX_TO_RAM_PIPELINE)
   ,.AXISTEN_IF_MSIX_FROM_RAM_PIPELINE(AXISTEN_IF_MSIX_FROM_RAM_PIPELINE)
   ,.AXISTEN_IF_MSIX_RX_PARITY_EN(AXISTEN_IF_MSIX_RX_PARITY_EN)
   ,.AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE(AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE)
   ,.AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT(AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT)
   ,.AXISTEN_IF_CQ_EN_POISONED_MEM_WR(AXISTEN_IF_CQ_EN_POISONED_MEM_WR)
   ,.PM_ASPML0S_TIMEOUT(PM_ASPML0S_TIMEOUT)
   ,.PM_L1_REENTRY_DELAY(PM_L1_REENTRY_DELAY)
   ,.PM_ASPML1_ENTRY_DELAY(PM_ASPML1_ENTRY_DELAY)
   ,.PM_ENABLE_SLOT_POWER_CAPTURE(PM_ENABLE_SLOT_POWER_CAPTURE)
   ,.PM_PME_SERVICE_TIMEOUT_DELAY(PM_PME_SERVICE_TIMEOUT_DELAY)
   ,.PM_PME_TURNOFF_ACK_DELAY(PM_PME_TURNOFF_ACK_DELAY)
   ,.PL_UPSTREAM_FACING(PL_UPSTREAM_FACING)
   ,.PL_LINK_CAP_MAX_LINK_WIDTH(PL_LINK_CAP_MAX_LINK_WIDTH)
   ,.PL_LINK_CAP_MAX_LINK_SPEED(PL_LINK_CAP_MAX_LINK_SPEED)
   ,.PL_DISABLE_DC_BALANCE(PL_DISABLE_DC_BALANCE)
   ,.PL_DISABLE_EI_INFER_IN_L0(PL_DISABLE_EI_INFER_IN_L0)
   ,.PL_N_FTS(PL_N_FTS)
   ,.PL_DISABLE_UPCONFIG_CAPABLE(PL_DISABLE_UPCONFIG_CAPABLE)
   ,.PL_DISABLE_RETRAIN_ON_FRAMING_ERROR(PL_DISABLE_RETRAIN_ON_FRAMING_ERROR)
   ,.PL_DISABLE_RETRAIN_ON_EB_ERROR(PL_DISABLE_RETRAIN_ON_EB_ERROR)
   ,.PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR(PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR)
   ,.PL_REPORT_ALL_PHY_ERRORS(PL_REPORT_ALL_PHY_ERRORS)
   ,.PL_DISABLE_LFSR_UPDATE_ON_SKP(PL_DISABLE_LFSR_UPDATE_ON_SKP)
   ,.PL_LANE0_EQ_CONTROL(PL_LANE0_EQ_CONTROL)
   ,.PL_LANE1_EQ_CONTROL(PL_LANE1_EQ_CONTROL)
   ,.PL_LANE2_EQ_CONTROL(PL_LANE2_EQ_CONTROL)
   ,.PL_LANE3_EQ_CONTROL(PL_LANE3_EQ_CONTROL)
   ,.PL_LANE4_EQ_CONTROL(PL_LANE4_EQ_CONTROL)
   ,.PL_LANE5_EQ_CONTROL(PL_LANE5_EQ_CONTROL)
   ,.PL_LANE6_EQ_CONTROL(PL_LANE6_EQ_CONTROL)
   ,.PL_LANE7_EQ_CONTROL(PL_LANE7_EQ_CONTROL)
   ,.PL_LANE8_EQ_CONTROL(PL_LANE8_EQ_CONTROL)
   ,.PL_LANE9_EQ_CONTROL(PL_LANE9_EQ_CONTROL)
   ,.PL_LANE10_EQ_CONTROL(PL_LANE10_EQ_CONTROL)
   ,.PL_LANE11_EQ_CONTROL(PL_LANE11_EQ_CONTROL)
   ,.PL_LANE12_EQ_CONTROL(PL_LANE12_EQ_CONTROL)
   ,.PL_LANE13_EQ_CONTROL(PL_LANE13_EQ_CONTROL)
   ,.PL_LANE14_EQ_CONTROL(PL_LANE14_EQ_CONTROL)
   ,.PL_LANE15_EQ_CONTROL(PL_LANE15_EQ_CONTROL)
   ,.PL_EQ_BYPASS_PHASE23(PL_EQ_BYPASS_PHASE23)
   ,.PL_EQ_ADAPT_ITER_COUNT(PL_EQ_ADAPT_ITER_COUNT)
   ,.PL_EQ_ADAPT_REJECT_RETRY_COUNT(PL_EQ_ADAPT_REJECT_RETRY_COUNT)
   ,.PL_EQ_SHORT_ADAPT_PHASE(PL_EQ_SHORT_ADAPT_PHASE)
   ,.PL_EQ_ADAPT_DISABLE_COEFF_CHECK(PL_EQ_ADAPT_DISABLE_COEFF_CHECK)
   ,.PL_EQ_ADAPT_DISABLE_PRESET_CHECK(PL_EQ_ADAPT_DISABLE_PRESET_CHECK)
   ,.PL_EQ_DEFAULT_TX_PRESET(PL_EQ_DEFAULT_TX_PRESET)
   ,.PL_EQ_DEFAULT_RX_PRESET_HINT(PL_EQ_DEFAULT_RX_PRESET_HINT)
   ,.PL_EQ_RX_ADAPT_EQ_PHASE0(PL_EQ_RX_ADAPT_EQ_PHASE0)
   ,.PL_EQ_RX_ADAPT_EQ_PHASE1(PL_EQ_RX_ADAPT_EQ_PHASE1)
   ,.PL_EQ_DISABLE_MISMATCH_CHECK(PL_EQ_DISABLE_MISMATCH_CHECK)
   ,.PL_RX_L0S_EXIT_TO_RECOVERY(PL_RX_L0S_EXIT_TO_RECOVERY)
   ,.PL_EQ_TX_8G_EQ_TS2_ENABLE(PL_EQ_TX_8G_EQ_TS2_ENABLE)
   ,.PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4(PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4)
   ,.PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3(PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3)
   ,.PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2(PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2)
   ,.PL_DESKEW_ON_SKIP_IN_GEN12(PL_DESKEW_ON_SKIP_IN_GEN12)
   ,.PL_INFER_EI_DISABLE_REC_RC(PL_INFER_EI_DISABLE_REC_RC)
   ,.PL_INFER_EI_DISABLE_REC_SPD(PL_INFER_EI_DISABLE_REC_SPD)
   ,.PL_INFER_EI_DISABLE_LPBK_ACTIVE(PL_INFER_EI_DISABLE_LPBK_ACTIVE)
   ,.PL_RX_ADAPT_TIMER_RRL_GEN3(PL_RX_ADAPT_TIMER_RRL_GEN3)
   ,.PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS(PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS)
   ,.PL_RX_ADAPT_TIMER_RRL_GEN4(PL_RX_ADAPT_TIMER_RRL_GEN4)
   ,.PL_RX_ADAPT_TIMER_CLWS_GEN3(PL_RX_ADAPT_TIMER_CLWS_GEN3)
   ,.PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS(PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS)
   ,.PL_RX_ADAPT_TIMER_CLWS_GEN4(PL_RX_ADAPT_TIMER_CLWS_GEN4)
   ,.PL_DISABLE_LANE_REVERSAL(PL_DISABLE_LANE_REVERSAL)
   ,.PL_CFG_STATE_ROBUSTNESS_ENABLE(PL_CFG_STATE_ROBUSTNESS_ENABLE)
   ,.PL_REDO_EQ_SOURCE_SELECT(PL_REDO_EQ_SOURCE_SELECT)
   ,.PL_DEEMPH_SOURCE_SELECT(PL_DEEMPH_SOURCE_SELECT)
   ,.PL_EXIT_LOOPBACK_ON_EI_ENTRY(PL_EXIT_LOOPBACK_ON_EI_ENTRY)
   ,.PL_QUIESCE_GUARANTEE_DISABLE(PL_QUIESCE_GUARANTEE_DISABLE)
   ,.PL_SRIS_ENABLE(PL_SRIS_ENABLE)
   ,.PL_SRIS_SKPOS_GEN_SPD_VEC(PL_SRIS_SKPOS_GEN_SPD_VEC)
   ,.PL_SRIS_SKPOS_REC_SPD_VEC(PL_SRIS_SKPOS_REC_SPD_VEC)
   ,.PL_SIM_FAST_LINK_TRAINING(PL_SIM_FAST_LINK_TRAINING)
   ,.PL_USER_SPARE(PL_USER_SPARE)
   ,.LL_ACK_TIMEOUT_EN(LL_ACK_TIMEOUT_EN)
   ,.LL_ACK_TIMEOUT(LL_ACK_TIMEOUT)
   ,.LL_ACK_TIMEOUT_FUNC(LL_ACK_TIMEOUT_FUNC)
   ,.LL_REPLAY_TIMEOUT_EN(LL_REPLAY_TIMEOUT_EN)
   ,.LL_REPLAY_TIMEOUT(LL_REPLAY_TIMEOUT)
   ,.LL_REPLAY_TIMEOUT_FUNC(LL_REPLAY_TIMEOUT_FUNC)
   ,.LL_REPLAY_TO_RAM_PIPELINE(LL_REPLAY_TO_RAM_PIPELINE)
   ,.LL_REPLAY_FROM_RAM_PIPELINE(LL_REPLAY_FROM_RAM_PIPELINE)
   ,.LL_DISABLE_SCHED_TX_NAK(LL_DISABLE_SCHED_TX_NAK)
   ,.LL_TX_TLP_PARITY_CHK(LL_TX_TLP_PARITY_CHK)
   ,.LL_RX_TLP_PARITY_GEN(LL_RX_TLP_PARITY_GEN)
   ,.LL_USER_SPARE(LL_USER_SPARE)
   ,.IS_SWITCH_PORT(IS_SWITCH_PORT)
   ,.CFG_BYPASS_MODE_ENABLE(CFG_BYPASS_MODE_ENABLE)
   ,.TL_PF_ENABLE_REG(TL_PF_ENABLE_REG)
   ,.TL_CREDITS_CD(TL_CREDITS_CD)
   ,.TL_CREDITS_CH(TL_CREDITS_CH)
   ,.TL_COMPLETION_RAM_SIZE(TL_COMPLETION_RAM_SIZE)
   ,.TL_COMPLETION_RAM_NUM_TLPS(TL_COMPLETION_RAM_NUM_TLPS)
   ,.TL_CREDITS_NPD(TL_CREDITS_NPD)
   ,.TL_CREDITS_NPH(TL_CREDITS_NPH)
   ,.TL_CREDITS_PD(TL_CREDITS_PD)
   ,.TL_CREDITS_PH(TL_CREDITS_PH)
   ,.TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE(TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE)
   ,.TL_RX_COMPLETION_TO_RAM_READ_PIPELINE(TL_RX_COMPLETION_TO_RAM_READ_PIPELINE)
   ,.TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE(TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE)
   ,.TL_POSTED_RAM_SIZE(TL_POSTED_RAM_SIZE)
   ,.TL_RX_POSTED_TO_RAM_WRITE_PIPELINE(TL_RX_POSTED_TO_RAM_WRITE_PIPELINE)
   ,.TL_RX_POSTED_TO_RAM_READ_PIPELINE(TL_RX_POSTED_TO_RAM_READ_PIPELINE)
   ,.TL_RX_POSTED_FROM_RAM_READ_PIPELINE(TL_RX_POSTED_FROM_RAM_READ_PIPELINE)
   ,.TL_TX_MUX_STRICT_PRIORITY(TL_TX_MUX_STRICT_PRIORITY)
   ,.TL_TX_TLP_STRADDLE_ENABLE(TL_TX_TLP_STRADDLE_ENABLE)
   ,.TL_TX_TLP_TERMINATE_PARITY(TL_TX_TLP_TERMINATE_PARITY)
   ,.TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT(TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT)
   ,.TL_FC_UPDATE_MIN_INTERVAL_TIME(TL_FC_UPDATE_MIN_INTERVAL_TIME)
   ,.TL_USER_SPARE(TL_USER_SPARE)
   ,.PF0_CLASS_CODE(PF0_CLASS_CODE)
   ,.PF1_CLASS_CODE(PF1_CLASS_CODE)
   ,.PF2_CLASS_CODE(PF2_CLASS_CODE)
   ,.PF3_CLASS_CODE(PF3_CLASS_CODE)
   ,.PF0_INTERRUPT_PIN(PF0_INTERRUPT_PIN)
   ,.PF1_INTERRUPT_PIN(PF1_INTERRUPT_PIN)
   ,.PF2_INTERRUPT_PIN(PF2_INTERRUPT_PIN)
   ,.PF3_INTERRUPT_PIN(PF3_INTERRUPT_PIN)
   ,.PF0_CAPABILITY_POINTER(PF0_CAPABILITY_POINTER)
   ,.PF1_CAPABILITY_POINTER(PF1_CAPABILITY_POINTER)
   ,.PF2_CAPABILITY_POINTER(PF2_CAPABILITY_POINTER)
   ,.PF3_CAPABILITY_POINTER(PF3_CAPABILITY_POINTER)
   ,.VF0_CAPABILITY_POINTER(VF0_CAPABILITY_POINTER)
   ,.LEGACY_CFG_EXTEND_INTERFACE_ENABLE(LEGACY_CFG_EXTEND_INTERFACE_ENABLE)
   ,.EXTENDED_CFG_EXTEND_INTERFACE_ENABLE(EXTENDED_CFG_EXTEND_INTERFACE_ENABLE)
   ,.TL2CFG_IF_PARITY_CHK(TL2CFG_IF_PARITY_CHK)
   ,.PF0_BAR0_CONTROL(PF0_BAR0_CONTROL)
   ,.PF1_BAR0_CONTROL(PF1_BAR0_CONTROL)
   ,.PF2_BAR0_CONTROL(PF2_BAR0_CONTROL)
   ,.PF3_BAR0_CONTROL(PF3_BAR0_CONTROL)
   ,.PF0_BAR0_APERTURE_SIZE(PF0_BAR0_APERTURE_SIZE)
   ,.PF1_BAR0_APERTURE_SIZE(PF1_BAR0_APERTURE_SIZE)
   ,.PF2_BAR0_APERTURE_SIZE(PF2_BAR0_APERTURE_SIZE)
   ,.PF3_BAR0_APERTURE_SIZE(PF3_BAR0_APERTURE_SIZE)
   ,.PF0_BAR1_CONTROL(PF0_BAR1_CONTROL)
   ,.PF1_BAR1_CONTROL(PF1_BAR1_CONTROL)
   ,.PF2_BAR1_CONTROL(PF2_BAR1_CONTROL)
   ,.PF3_BAR1_CONTROL(PF3_BAR1_CONTROL)
   ,.PF0_BAR1_APERTURE_SIZE(PF0_BAR1_APERTURE_SIZE)
   ,.PF1_BAR1_APERTURE_SIZE(PF1_BAR1_APERTURE_SIZE)
   ,.PF2_BAR1_APERTURE_SIZE(PF2_BAR1_APERTURE_SIZE)
   ,.PF3_BAR1_APERTURE_SIZE(PF3_BAR1_APERTURE_SIZE)
   ,.PF0_BAR2_CONTROL(PF0_BAR2_CONTROL)
   ,.PF1_BAR2_CONTROL(PF1_BAR2_CONTROL)
   ,.PF2_BAR2_CONTROL(PF2_BAR2_CONTROL)
   ,.PF3_BAR2_CONTROL(PF3_BAR2_CONTROL)
   ,.PF0_BAR2_APERTURE_SIZE(PF0_BAR2_APERTURE_SIZE)
   ,.PF1_BAR2_APERTURE_SIZE(PF1_BAR2_APERTURE_SIZE)
   ,.PF2_BAR2_APERTURE_SIZE(PF2_BAR2_APERTURE_SIZE)
   ,.PF3_BAR2_APERTURE_SIZE(PF3_BAR2_APERTURE_SIZE)
   ,.PF0_BAR3_CONTROL(PF0_BAR3_CONTROL)
   ,.PF1_BAR3_CONTROL(PF1_BAR3_CONTROL)
   ,.PF2_BAR3_CONTROL(PF2_BAR3_CONTROL)
   ,.PF3_BAR3_CONTROL(PF3_BAR3_CONTROL)
   ,.PF0_BAR3_APERTURE_SIZE(PF0_BAR3_APERTURE_SIZE)
   ,.PF1_BAR3_APERTURE_SIZE(PF1_BAR3_APERTURE_SIZE)
   ,.PF2_BAR3_APERTURE_SIZE(PF2_BAR3_APERTURE_SIZE)
   ,.PF3_BAR3_APERTURE_SIZE(PF3_BAR3_APERTURE_SIZE)
   ,.PF0_BAR4_CONTROL(PF0_BAR4_CONTROL)
   ,.PF1_BAR4_CONTROL(PF1_BAR4_CONTROL)
   ,.PF2_BAR4_CONTROL(PF2_BAR4_CONTROL)
   ,.PF3_BAR4_CONTROL(PF3_BAR4_CONTROL)
   ,.PF0_BAR4_APERTURE_SIZE(PF0_BAR4_APERTURE_SIZE)
   ,.PF1_BAR4_APERTURE_SIZE(PF1_BAR4_APERTURE_SIZE)
   ,.PF2_BAR4_APERTURE_SIZE(PF2_BAR4_APERTURE_SIZE)
   ,.PF3_BAR4_APERTURE_SIZE(PF3_BAR4_APERTURE_SIZE)
   ,.PF0_BAR5_CONTROL(PF0_BAR5_CONTROL)
   ,.PF1_BAR5_CONTROL(PF1_BAR5_CONTROL)
   ,.PF2_BAR5_CONTROL(PF2_BAR5_CONTROL)
   ,.PF3_BAR5_CONTROL(PF3_BAR5_CONTROL)
   ,.PF0_BAR5_APERTURE_SIZE(PF0_BAR5_APERTURE_SIZE)
   ,.PF1_BAR5_APERTURE_SIZE(PF1_BAR5_APERTURE_SIZE)
   ,.PF2_BAR5_APERTURE_SIZE(PF2_BAR5_APERTURE_SIZE)
   ,.PF3_BAR5_APERTURE_SIZE(PF3_BAR5_APERTURE_SIZE)
   ,.PF0_EXPANSION_ROM_ENABLE(PF0_EXPANSION_ROM_ENABLE)
   ,.PF1_EXPANSION_ROM_ENABLE(PF1_EXPANSION_ROM_ENABLE)
   ,.PF2_EXPANSION_ROM_ENABLE(PF2_EXPANSION_ROM_ENABLE)
   ,.PF3_EXPANSION_ROM_ENABLE(PF3_EXPANSION_ROM_ENABLE)
   ,.PF0_EXPANSION_ROM_APERTURE_SIZE(PF0_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF1_EXPANSION_ROM_APERTURE_SIZE(PF1_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF2_EXPANSION_ROM_APERTURE_SIZE(PF2_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF3_EXPANSION_ROM_APERTURE_SIZE(PF3_EXPANSION_ROM_APERTURE_SIZE)
   ,.PF0_PCIE_CAP_NEXTPTR(PF0_PCIE_CAP_NEXTPTR)
   ,.PF1_PCIE_CAP_NEXTPTR(PF1_PCIE_CAP_NEXTPTR)
   ,.PF2_PCIE_CAP_NEXTPTR(PF2_PCIE_CAP_NEXTPTR)
   ,.PF3_PCIE_CAP_NEXTPTR(PF3_PCIE_CAP_NEXTPTR)
   ,.VFG0_PCIE_CAP_NEXTPTR(VFG0_PCIE_CAP_NEXTPTR)
   ,.VFG1_PCIE_CAP_NEXTPTR(VFG1_PCIE_CAP_NEXTPTR)
   ,.VFG2_PCIE_CAP_NEXTPTR(VFG2_PCIE_CAP_NEXTPTR)
   ,.VFG3_PCIE_CAP_NEXTPTR(VFG3_PCIE_CAP_NEXTPTR)
   ,.HEADER_TYPE_OVERRIDE(HEADER_TYPE_OVERRIDE)
   ,.PF0_LINK_CONTROL_RCB(PF0_LINK_CONTROL_RCB)
   ,.PF0_DEV_CAP_MAX_PAYLOAD_SIZE(PF0_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF1_DEV_CAP_MAX_PAYLOAD_SIZE(PF1_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF2_DEV_CAP_MAX_PAYLOAD_SIZE(PF2_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF3_DEV_CAP_MAX_PAYLOAD_SIZE(PF3_DEV_CAP_MAX_PAYLOAD_SIZE)
   ,.PF0_DEV_CAP_EXT_TAG_SUPPORTED(PF0_DEV_CAP_EXT_TAG_SUPPORTED)
   ,.PF0_DEV_CAP_ENDPOINT_L0S_LATENCY(PF0_DEV_CAP_ENDPOINT_L0S_LATENCY)
   ,.PF0_DEV_CAP_ENDPOINT_L1_LATENCY(PF0_DEV_CAP_ENDPOINT_L1_LATENCY)
   ,.PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE(PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE)
   ,.PF0_LINK_CAP_ASPM_SUPPORT(PF0_LINK_CAP_ASPM_SUPPORT)
   ,.PF0_LINK_STATUS_SLOT_CLOCK_CONFIG(PF0_LINK_STATUS_SLOT_CLOCK_CONFIG)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4(PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3)
   ,.PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4(PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4(PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3)
   ,.PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4(PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4)
   ,.PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE(PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE)
   ,.PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT(PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT(PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT(PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_LTR_SUPPORT(PF0_DEV_CAP2_LTR_SUPPORT)
   ,.PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT(PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT)
   ,.PF0_DEV_CAP2_OBFF_SUPPORT(PF0_DEV_CAP2_OBFF_SUPPORT)
   ,.PF0_DEV_CAP2_ARI_FORWARD_ENABLE(PF0_DEV_CAP2_ARI_FORWARD_ENABLE)
   ,.PF0_MSI_CAP_NEXTPTR(PF0_MSI_CAP_NEXTPTR)
   ,.PF1_MSI_CAP_NEXTPTR(PF1_MSI_CAP_NEXTPTR)
   ,.PF2_MSI_CAP_NEXTPTR(PF2_MSI_CAP_NEXTPTR)
   ,.PF3_MSI_CAP_NEXTPTR(PF3_MSI_CAP_NEXTPTR)
   ,.PF0_MSI_CAP_PERVECMASKCAP(PF0_MSI_CAP_PERVECMASKCAP)
   ,.PF1_MSI_CAP_PERVECMASKCAP(PF1_MSI_CAP_PERVECMASKCAP)
   ,.PF2_MSI_CAP_PERVECMASKCAP(PF2_MSI_CAP_PERVECMASKCAP)
   ,.PF3_MSI_CAP_PERVECMASKCAP(PF3_MSI_CAP_PERVECMASKCAP)
   ,.PF0_MSI_CAP_MULTIMSGCAP(PF0_MSI_CAP_MULTIMSGCAP)
   ,.PF1_MSI_CAP_MULTIMSGCAP(PF1_MSI_CAP_MULTIMSGCAP)
   ,.PF2_MSI_CAP_MULTIMSGCAP(PF2_MSI_CAP_MULTIMSGCAP)
   ,.PF3_MSI_CAP_MULTIMSGCAP(PF3_MSI_CAP_MULTIMSGCAP)
   ,.PF0_MSIX_CAP_NEXTPTR(PF0_MSIX_CAP_NEXTPTR)
   ,.PF1_MSIX_CAP_NEXTPTR(PF1_MSIX_CAP_NEXTPTR)
   ,.PF2_MSIX_CAP_NEXTPTR(PF2_MSIX_CAP_NEXTPTR)
   ,.PF3_MSIX_CAP_NEXTPTR(PF3_MSIX_CAP_NEXTPTR)
   ,.VFG0_MSIX_CAP_NEXTPTR(VFG0_MSIX_CAP_NEXTPTR)
   ,.VFG1_MSIX_CAP_NEXTPTR(VFG1_MSIX_CAP_NEXTPTR)
   ,.VFG2_MSIX_CAP_NEXTPTR(VFG2_MSIX_CAP_NEXTPTR)
   ,.VFG3_MSIX_CAP_NEXTPTR(VFG3_MSIX_CAP_NEXTPTR)
   ,.PF0_MSIX_CAP_PBA_BIR(PF0_MSIX_CAP_PBA_BIR)
   ,.PF1_MSIX_CAP_PBA_BIR(PF1_MSIX_CAP_PBA_BIR)
   ,.PF2_MSIX_CAP_PBA_BIR(PF2_MSIX_CAP_PBA_BIR)
   ,.PF3_MSIX_CAP_PBA_BIR(PF3_MSIX_CAP_PBA_BIR)
   ,.VFG0_MSIX_CAP_PBA_BIR(VFG0_MSIX_CAP_PBA_BIR)
   ,.VFG1_MSIX_CAP_PBA_BIR(VFG1_MSIX_CAP_PBA_BIR)
   ,.VFG2_MSIX_CAP_PBA_BIR(VFG2_MSIX_CAP_PBA_BIR)
   ,.VFG3_MSIX_CAP_PBA_BIR(VFG3_MSIX_CAP_PBA_BIR)
   ,.PF0_MSIX_CAP_PBA_OFFSET(PF0_MSIX_CAP_PBA_OFFSET)
   ,.PF1_MSIX_CAP_PBA_OFFSET(PF1_MSIX_CAP_PBA_OFFSET)
   ,.PF2_MSIX_CAP_PBA_OFFSET(PF2_MSIX_CAP_PBA_OFFSET)
   ,.PF3_MSIX_CAP_PBA_OFFSET(PF3_MSIX_CAP_PBA_OFFSET)
   ,.VFG0_MSIX_CAP_PBA_OFFSET(VFG0_MSIX_CAP_PBA_OFFSET)
   ,.VFG1_MSIX_CAP_PBA_OFFSET(VFG1_MSIX_CAP_PBA_OFFSET)
   ,.VFG2_MSIX_CAP_PBA_OFFSET(VFG2_MSIX_CAP_PBA_OFFSET)
   ,.VFG3_MSIX_CAP_PBA_OFFSET(VFG3_MSIX_CAP_PBA_OFFSET)
   ,.PF0_MSIX_CAP_TABLE_BIR(PF0_MSIX_CAP_TABLE_BIR)
   ,.PF1_MSIX_CAP_TABLE_BIR(PF1_MSIX_CAP_TABLE_BIR)
   ,.PF2_MSIX_CAP_TABLE_BIR(PF2_MSIX_CAP_TABLE_BIR)
   ,.PF3_MSIX_CAP_TABLE_BIR(PF3_MSIX_CAP_TABLE_BIR)
   ,.VFG0_MSIX_CAP_TABLE_BIR(VFG0_MSIX_CAP_TABLE_BIR)
   ,.VFG1_MSIX_CAP_TABLE_BIR(VFG1_MSIX_CAP_TABLE_BIR)
   ,.VFG2_MSIX_CAP_TABLE_BIR(VFG2_MSIX_CAP_TABLE_BIR)
   ,.VFG3_MSIX_CAP_TABLE_BIR(VFG3_MSIX_CAP_TABLE_BIR)
   ,.PF0_MSIX_CAP_TABLE_OFFSET(PF0_MSIX_CAP_TABLE_OFFSET)
   ,.PF1_MSIX_CAP_TABLE_OFFSET(PF1_MSIX_CAP_TABLE_OFFSET)
   ,.PF2_MSIX_CAP_TABLE_OFFSET(PF2_MSIX_CAP_TABLE_OFFSET)
   ,.PF3_MSIX_CAP_TABLE_OFFSET(PF3_MSIX_CAP_TABLE_OFFSET)
   ,.VFG0_MSIX_CAP_TABLE_OFFSET(VFG0_MSIX_CAP_TABLE_OFFSET)
   ,.VFG1_MSIX_CAP_TABLE_OFFSET(VFG1_MSIX_CAP_TABLE_OFFSET)
   ,.VFG2_MSIX_CAP_TABLE_OFFSET(VFG2_MSIX_CAP_TABLE_OFFSET)
   ,.VFG3_MSIX_CAP_TABLE_OFFSET(VFG3_MSIX_CAP_TABLE_OFFSET)
   ,.PF0_MSIX_CAP_TABLE_SIZE(PF0_MSIX_CAP_TABLE_SIZE)
   ,.PF1_MSIX_CAP_TABLE_SIZE(PF1_MSIX_CAP_TABLE_SIZE)
   ,.PF2_MSIX_CAP_TABLE_SIZE(PF2_MSIX_CAP_TABLE_SIZE)
   ,.PF3_MSIX_CAP_TABLE_SIZE(PF3_MSIX_CAP_TABLE_SIZE)
   ,.VFG0_MSIX_CAP_TABLE_SIZE(VFG0_MSIX_CAP_TABLE_SIZE)
   ,.VFG1_MSIX_CAP_TABLE_SIZE(VFG1_MSIX_CAP_TABLE_SIZE)
   ,.VFG2_MSIX_CAP_TABLE_SIZE(VFG2_MSIX_CAP_TABLE_SIZE)
   ,.VFG3_MSIX_CAP_TABLE_SIZE(VFG3_MSIX_CAP_TABLE_SIZE)
   ,.PF0_MSIX_VECTOR_COUNT(PF0_MSIX_VECTOR_COUNT)
   ,.PF0_PM_CAP_ID(PF0_PM_CAP_ID)
   ,.PF0_PM_CAP_NEXTPTR(PF0_PM_CAP_NEXTPTR)
   ,.PF1_PM_CAP_NEXTPTR(PF1_PM_CAP_NEXTPTR)
   ,.PF2_PM_CAP_NEXTPTR(PF2_PM_CAP_NEXTPTR)
   ,.PF3_PM_CAP_NEXTPTR(PF3_PM_CAP_NEXTPTR)
   ,.PF0_PM_CAP_PMESUPPORT_D3HOT(PF0_PM_CAP_PMESUPPORT_D3HOT)
   ,.PF0_PM_CAP_PMESUPPORT_D1(PF0_PM_CAP_PMESUPPORT_D1)
   ,.PF0_PM_CAP_PMESUPPORT_D0(PF0_PM_CAP_PMESUPPORT_D0)
   ,.PF0_PM_CAP_SUPP_D1_STATE(PF0_PM_CAP_SUPP_D1_STATE)
   ,.PF0_PM_CAP_VER_ID(PF0_PM_CAP_VER_ID)
   ,.PF0_PM_CSR_NOSOFTRESET(PF0_PM_CSR_NOSOFTRESET)
   ,.PM_ENABLE_L23_ENTRY(PM_ENABLE_L23_ENTRY)
   ,.DNSTREAM_LINK_NUM(DNSTREAM_LINK_NUM)
   ,.AUTO_FLR_RESPONSE(AUTO_FLR_RESPONSE)
   ,.PF0_DSN_CAP_NEXTPTR(PF0_DSN_CAP_NEXTPTR)
   ,.PF1_DSN_CAP_NEXTPTR(PF1_DSN_CAP_NEXTPTR)
   ,.PF2_DSN_CAP_NEXTPTR(PF2_DSN_CAP_NEXTPTR)
   ,.PF3_DSN_CAP_NEXTPTR(PF3_DSN_CAP_NEXTPTR)
   ,.DSN_CAP_ENABLE(DSN_CAP_ENABLE)
   ,.PF0_VC_CAP_VER(PF0_VC_CAP_VER)
   ,.PF0_VC_CAP_NEXTPTR(PF0_VC_CAP_NEXTPTR)
   ,.PF0_VC_CAP_ENABLE(PF0_VC_CAP_ENABLE)
   ,.PF0_SECONDARY_PCIE_CAP_NEXTPTR(PF0_SECONDARY_PCIE_CAP_NEXTPTR)
   ,.PF0_AER_CAP_NEXTPTR(PF0_AER_CAP_NEXTPTR)
   ,.PF1_AER_CAP_NEXTPTR(PF1_AER_CAP_NEXTPTR)
   ,.PF2_AER_CAP_NEXTPTR(PF2_AER_CAP_NEXTPTR)
   ,.PF3_AER_CAP_NEXTPTR(PF3_AER_CAP_NEXTPTR)
   ,.PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE(PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE)
   ,.ARI_CAP_ENABLE(ARI_CAP_ENABLE)
   ,.PF0_ARI_CAP_NEXTPTR(PF0_ARI_CAP_NEXTPTR)
   ,.PF1_ARI_CAP_NEXTPTR(PF1_ARI_CAP_NEXTPTR)
   ,.PF2_ARI_CAP_NEXTPTR(PF2_ARI_CAP_NEXTPTR)
   ,.PF3_ARI_CAP_NEXTPTR(PF3_ARI_CAP_NEXTPTR)
   ,.VFG0_ARI_CAP_NEXTPTR(VFG0_ARI_CAP_NEXTPTR)
   ,.VFG1_ARI_CAP_NEXTPTR(VFG1_ARI_CAP_NEXTPTR)
   ,.VFG2_ARI_CAP_NEXTPTR(VFG2_ARI_CAP_NEXTPTR)
   ,.VFG3_ARI_CAP_NEXTPTR(VFG3_ARI_CAP_NEXTPTR)
   ,.PF0_ARI_CAP_VER(PF0_ARI_CAP_VER)
   ,.PF0_ARI_CAP_NEXT_FUNC(PF0_ARI_CAP_NEXT_FUNC)
   ,.PF1_ARI_CAP_NEXT_FUNC(PF1_ARI_CAP_NEXT_FUNC)
   ,.PF2_ARI_CAP_NEXT_FUNC(PF2_ARI_CAP_NEXT_FUNC)
   ,.PF3_ARI_CAP_NEXT_FUNC(PF3_ARI_CAP_NEXT_FUNC)
   ,.PF0_LTR_CAP_NEXTPTR(PF0_LTR_CAP_NEXTPTR)
   ,.PF0_LTR_CAP_VER(PF0_LTR_CAP_VER)
   ,.PF0_LTR_CAP_MAX_SNOOP_LAT(PF0_LTR_CAP_MAX_SNOOP_LAT)
   ,.PF0_LTR_CAP_MAX_NOSNOOP_LAT(PF0_LTR_CAP_MAX_NOSNOOP_LAT)
   ,.LTR_TX_MESSAGE_ON_LTR_ENABLE(LTR_TX_MESSAGE_ON_LTR_ENABLE)
   ,.LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE(LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE)
   ,.LTR_TX_MESSAGE_MINIMUM_INTERVAL(LTR_TX_MESSAGE_MINIMUM_INTERVAL)
   ,.SRIOV_CAP_ENABLE(SRIOV_CAP_ENABLE)
   ,.PF0_SRIOV_CAP_NEXTPTR(PF0_SRIOV_CAP_NEXTPTR)
   ,.PF1_SRIOV_CAP_NEXTPTR(PF1_SRIOV_CAP_NEXTPTR)
   ,.PF2_SRIOV_CAP_NEXTPTR(PF2_SRIOV_CAP_NEXTPTR)
   ,.PF3_SRIOV_CAP_NEXTPTR(PF3_SRIOV_CAP_NEXTPTR)
   ,.PF0_SRIOV_CAP_VER(PF0_SRIOV_CAP_VER)
   ,.PF1_SRIOV_CAP_VER(PF1_SRIOV_CAP_VER)
   ,.PF2_SRIOV_CAP_VER(PF2_SRIOV_CAP_VER)
   ,.PF3_SRIOV_CAP_VER(PF3_SRIOV_CAP_VER)
   ,.PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED(PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED)
   ,.PF0_SRIOV_CAP_INITIAL_VF(PF0_SRIOV_CAP_INITIAL_VF)
   ,.PF1_SRIOV_CAP_INITIAL_VF(PF1_SRIOV_CAP_INITIAL_VF)
   ,.PF2_SRIOV_CAP_INITIAL_VF(PF2_SRIOV_CAP_INITIAL_VF)
   ,.PF3_SRIOV_CAP_INITIAL_VF(PF3_SRIOV_CAP_INITIAL_VF)
   ,.PF0_SRIOV_CAP_TOTAL_VF(PF0_SRIOV_CAP_TOTAL_VF)
   ,.PF1_SRIOV_CAP_TOTAL_VF(PF1_SRIOV_CAP_TOTAL_VF)
   ,.PF2_SRIOV_CAP_TOTAL_VF(PF2_SRIOV_CAP_TOTAL_VF)
   ,.PF3_SRIOV_CAP_TOTAL_VF(PF3_SRIOV_CAP_TOTAL_VF)
   ,.PF0_SRIOV_FUNC_DEP_LINK(PF0_SRIOV_FUNC_DEP_LINK)
   ,.PF1_SRIOV_FUNC_DEP_LINK(PF1_SRIOV_FUNC_DEP_LINK)
   ,.PF2_SRIOV_FUNC_DEP_LINK(PF2_SRIOV_FUNC_DEP_LINK)
   ,.PF3_SRIOV_FUNC_DEP_LINK(PF3_SRIOV_FUNC_DEP_LINK)
   ,.PF0_SRIOV_FIRST_VF_OFFSET(PF0_SRIOV_FIRST_VF_OFFSET)
   ,.PF1_SRIOV_FIRST_VF_OFFSET(PF1_SRIOV_FIRST_VF_OFFSET)
   ,.PF2_SRIOV_FIRST_VF_OFFSET(PF2_SRIOV_FIRST_VF_OFFSET)
   ,.PF3_SRIOV_FIRST_VF_OFFSET(PF3_SRIOV_FIRST_VF_OFFSET)
   ,.PF0_SRIOV_VF_DEVICE_ID(PF0_SRIOV_VF_DEVICE_ID)
   ,.PF1_SRIOV_VF_DEVICE_ID(PF1_SRIOV_VF_DEVICE_ID)
   ,.PF2_SRIOV_VF_DEVICE_ID(PF2_SRIOV_VF_DEVICE_ID)
   ,.PF3_SRIOV_VF_DEVICE_ID(PF3_SRIOV_VF_DEVICE_ID)
   ,.PF0_SRIOV_SUPPORTED_PAGE_SIZE(PF0_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF1_SRIOV_SUPPORTED_PAGE_SIZE(PF1_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF2_SRIOV_SUPPORTED_PAGE_SIZE(PF2_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF3_SRIOV_SUPPORTED_PAGE_SIZE(PF3_SRIOV_SUPPORTED_PAGE_SIZE)
   ,.PF0_SRIOV_BAR0_CONTROL(PF0_SRIOV_BAR0_CONTROL)
   ,.PF1_SRIOV_BAR0_CONTROL(PF1_SRIOV_BAR0_CONTROL)
   ,.PF2_SRIOV_BAR0_CONTROL(PF2_SRIOV_BAR0_CONTROL)
   ,.PF3_SRIOV_BAR0_CONTROL(PF3_SRIOV_BAR0_CONTROL)
   ,.PF0_SRIOV_BAR0_APERTURE_SIZE(PF0_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR0_APERTURE_SIZE(PF1_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR0_APERTURE_SIZE(PF2_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR0_APERTURE_SIZE(PF3_SRIOV_BAR0_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR1_CONTROL(PF0_SRIOV_BAR1_CONTROL)
   ,.PF1_SRIOV_BAR1_CONTROL(PF1_SRIOV_BAR1_CONTROL)
   ,.PF2_SRIOV_BAR1_CONTROL(PF2_SRIOV_BAR1_CONTROL)
   ,.PF3_SRIOV_BAR1_CONTROL(PF3_SRIOV_BAR1_CONTROL)
   ,.PF0_SRIOV_BAR1_APERTURE_SIZE(PF0_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR1_APERTURE_SIZE(PF1_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR1_APERTURE_SIZE(PF2_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR1_APERTURE_SIZE(PF3_SRIOV_BAR1_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR2_CONTROL(PF0_SRIOV_BAR2_CONTROL)
   ,.PF1_SRIOV_BAR2_CONTROL(PF1_SRIOV_BAR2_CONTROL)
   ,.PF2_SRIOV_BAR2_CONTROL(PF2_SRIOV_BAR2_CONTROL)
   ,.PF3_SRIOV_BAR2_CONTROL(PF3_SRIOV_BAR2_CONTROL)
   ,.PF0_SRIOV_BAR2_APERTURE_SIZE(PF0_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR2_APERTURE_SIZE(PF1_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR2_APERTURE_SIZE(PF2_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR2_APERTURE_SIZE(PF3_SRIOV_BAR2_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR3_CONTROL(PF0_SRIOV_BAR3_CONTROL)
   ,.PF1_SRIOV_BAR3_CONTROL(PF1_SRIOV_BAR3_CONTROL)
   ,.PF2_SRIOV_BAR3_CONTROL(PF2_SRIOV_BAR3_CONTROL)
   ,.PF3_SRIOV_BAR3_CONTROL(PF3_SRIOV_BAR3_CONTROL)
   ,.PF0_SRIOV_BAR3_APERTURE_SIZE(PF0_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR3_APERTURE_SIZE(PF1_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR3_APERTURE_SIZE(PF2_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR3_APERTURE_SIZE(PF3_SRIOV_BAR3_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR4_CONTROL(PF0_SRIOV_BAR4_CONTROL)
   ,.PF1_SRIOV_BAR4_CONTROL(PF1_SRIOV_BAR4_CONTROL)
   ,.PF2_SRIOV_BAR4_CONTROL(PF2_SRIOV_BAR4_CONTROL)
   ,.PF3_SRIOV_BAR4_CONTROL(PF3_SRIOV_BAR4_CONTROL)
   ,.PF0_SRIOV_BAR4_APERTURE_SIZE(PF0_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR4_APERTURE_SIZE(PF1_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR4_APERTURE_SIZE(PF2_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR4_APERTURE_SIZE(PF3_SRIOV_BAR4_APERTURE_SIZE)
   ,.PF0_SRIOV_BAR5_CONTROL(PF0_SRIOV_BAR5_CONTROL)
   ,.PF1_SRIOV_BAR5_CONTROL(PF1_SRIOV_BAR5_CONTROL)
   ,.PF2_SRIOV_BAR5_CONTROL(PF2_SRIOV_BAR5_CONTROL)
   ,.PF3_SRIOV_BAR5_CONTROL(PF3_SRIOV_BAR5_CONTROL)
   ,.PF0_SRIOV_BAR5_APERTURE_SIZE(PF0_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF1_SRIOV_BAR5_APERTURE_SIZE(PF1_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF2_SRIOV_BAR5_APERTURE_SIZE(PF2_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF3_SRIOV_BAR5_APERTURE_SIZE(PF3_SRIOV_BAR5_APERTURE_SIZE)
   ,.PF0_TPHR_CAP_NEXTPTR(PF0_TPHR_CAP_NEXTPTR)
   ,.PF1_TPHR_CAP_NEXTPTR(PF1_TPHR_CAP_NEXTPTR)
   ,.PF2_TPHR_CAP_NEXTPTR(PF2_TPHR_CAP_NEXTPTR)
   ,.PF3_TPHR_CAP_NEXTPTR(PF3_TPHR_CAP_NEXTPTR)
   ,.VFG0_TPHR_CAP_NEXTPTR(VFG0_TPHR_CAP_NEXTPTR)
   ,.VFG1_TPHR_CAP_NEXTPTR(VFG1_TPHR_CAP_NEXTPTR)
   ,.VFG2_TPHR_CAP_NEXTPTR(VFG2_TPHR_CAP_NEXTPTR)
   ,.VFG3_TPHR_CAP_NEXTPTR(VFG3_TPHR_CAP_NEXTPTR)
   ,.PF0_TPHR_CAP_VER(PF0_TPHR_CAP_VER)
   ,.PF0_TPHR_CAP_INT_VEC_MODE(PF0_TPHR_CAP_INT_VEC_MODE)
   ,.PF0_TPHR_CAP_DEV_SPECIFIC_MODE(PF0_TPHR_CAP_DEV_SPECIFIC_MODE)
   ,.PF0_TPHR_CAP_ST_TABLE_LOC(PF0_TPHR_CAP_ST_TABLE_LOC)
   ,.PF0_TPHR_CAP_ST_TABLE_SIZE(PF0_TPHR_CAP_ST_TABLE_SIZE)
   ,.PF0_TPHR_CAP_ST_MODE_SEL(PF0_TPHR_CAP_ST_MODE_SEL)
   ,.PF1_TPHR_CAP_ST_MODE_SEL(PF1_TPHR_CAP_ST_MODE_SEL)
   ,.PF2_TPHR_CAP_ST_MODE_SEL(PF2_TPHR_CAP_ST_MODE_SEL)
   ,.PF3_TPHR_CAP_ST_MODE_SEL(PF3_TPHR_CAP_ST_MODE_SEL)
   ,.VFG0_TPHR_CAP_ST_MODE_SEL(VFG0_TPHR_CAP_ST_MODE_SEL)
   ,.VFG1_TPHR_CAP_ST_MODE_SEL(VFG1_TPHR_CAP_ST_MODE_SEL)
   ,.VFG2_TPHR_CAP_ST_MODE_SEL(VFG2_TPHR_CAP_ST_MODE_SEL)
   ,.VFG3_TPHR_CAP_ST_MODE_SEL(VFG3_TPHR_CAP_ST_MODE_SEL)
   ,.PF0_TPHR_CAP_ENABLE(PF0_TPHR_CAP_ENABLE)
   ,.TPH_TO_RAM_PIPELINE(TPH_TO_RAM_PIPELINE)
   ,.TPH_FROM_RAM_PIPELINE(TPH_FROM_RAM_PIPELINE)
   ,.MCAP_ENABLE(MCAP_ENABLE)
   ,.MCAP_CONFIGURE_OVERRIDE(MCAP_CONFIGURE_OVERRIDE)
   ,.MCAP_CAP_NEXTPTR(MCAP_CAP_NEXTPTR)
   ,.MCAP_VSEC_ID(MCAP_VSEC_ID)
   ,.MCAP_VSEC_REV(MCAP_VSEC_REV)
   ,.MCAP_VSEC_LEN(MCAP_VSEC_LEN)
   ,.MCAP_FPGA_BITSTREAM_VERSION(MCAP_FPGA_BITSTREAM_VERSION)
   ,.MCAP_INTERRUPT_ON_MCAP_EOS(MCAP_INTERRUPT_ON_MCAP_EOS)
   ,.MCAP_INTERRUPT_ON_MCAP_ERROR(MCAP_INTERRUPT_ON_MCAP_ERROR)
   ,.MCAP_INPUT_GATE_DESIGN_SWITCH(MCAP_INPUT_GATE_DESIGN_SWITCH)
   ,.MCAP_EOS_DESIGN_SWITCH(MCAP_EOS_DESIGN_SWITCH)
   ,.MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH(MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH)
   ,.MCAP_GATE_IO_ENABLE_DESIGN_SWITCH(MCAP_GATE_IO_ENABLE_DESIGN_SWITCH)
   ,.SIM_JTAG_IDCODE(SIM_JTAG_IDCODE)
   ,.DEBUG_AXIST_DISABLE_FEATURE_BIT(DEBUG_AXIST_DISABLE_FEATURE_BIT)
   ,.DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS(DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS)
   ,.DEBUG_TL_DISABLE_FC_TIMEOUT(DEBUG_TL_DISABLE_FC_TIMEOUT)
   ,.DEBUG_PL_DISABLE_SCRAMBLING(DEBUG_PL_DISABLE_SCRAMBLING)
   ,.DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL (DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL )
   ,.DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW (DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW )
   ,.DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR(DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR)
   ,.DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR(DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR)
   ,.DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR(DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR)
   ,.DEBUG_PL_SIM_RESET_LFSR(DEBUG_PL_SIM_RESET_LFSR)
   ,.DEBUG_PL_SPARE(DEBUG_PL_SPARE)
   ,.DEBUG_LL_SPARE(DEBUG_LL_SPARE)
   ,.DEBUG_TL_SPARE(DEBUG_TL_SPARE)
   ,.DEBUG_AXI4ST_SPARE(DEBUG_AXI4ST_SPARE)
   ,.DEBUG_CFG_SPARE(DEBUG_CFG_SPARE)
   ,.DEBUG_CAR_SPARE(DEBUG_CAR_SPARE)
   ,.SPARE_BIT0(AXISTEN_IF_RQ_CC_REGISTERED_TREADY)
   ,.SPARE_BIT1(SPARE_BIT1)
   ,.SPARE_BIT2(SPARE_BIT2)
   ,.SPARE_BIT3(SPARE_BIT3)
   ,.SPARE_BIT4(SPARE_BIT4)
   ,.SPARE_BIT5(SPARE_BIT5)
   ,.SPARE_BIT6(SPARE_BIT6)
   ,.SPARE_BIT7(SPARE_BIT7)
   ,.SPARE_BIT8(SPARE_BIT8)
   ,.SPARE_BYTE0(SPARE_BYTE0)
   ,.SPARE_BYTE1(SPARE_BYTE1)
   ,.SPARE_BYTE2(SPARE_BYTE2)
   ,.SPARE_BYTE3(SPARE_BYTE3)
   ,.SPARE_WORD0(SPARE_WORD0)
   ,.SPARE_WORD1(SPARE_WORD1)
   ,.SPARE_WORD2(SPARE_WORD2)
   ,.SPARE_WORD3(SPARE_WORD3)

  ) pcie_4_0_e4_inst ( 

    .AXIUSERIN(axi_user_in[7:0])
   ,.AXIUSEROUT(axi_user_out[7:0])
   ,.CFGBUSNUMBER(cfg_bus_number[7:0])
   ,.CFGCONFIGSPACEENABLE(cfg_config_space_enable)
   ,.CFGCURRENTSPEED(cfg_current_speed[1:0])
   ,.CFGDEVIDPF0(cfg_dev_id_pf0[15:0])
   ,.CFGDEVIDPF1(cfg_dev_id_pf1[15:0])
   ,.CFGDEVIDPF2(cfg_dev_id_pf2[15:0])
   ,.CFGDEVIDPF3(cfg_dev_id_pf3[15:0])
   ,.CFGDSBUSNUMBER(cfg_ds_bus_number[7:0])
   ,.CFGDSDEVICENUMBER(cfg_ds_device_number[4:0])
   ,.CFGDSFUNCTIONNUMBER(cfg_ds_function_number[2:0])
   ,.CFGDSN(cfg_dsn[63:0])
   ,.CFGDSPORTNUMBER(cfg_ds_port_number[7:0])
   ,.CFGERRCORIN(cfg_err_cor_in)
   ,.CFGERRCOROUT(cfg_err_cor_out)
   ,.CFGERRFATALOUT(cfg_err_fatal_out)
   ,.CFGERRNONFATALOUT(cfg_err_nonfatal_out)
   ,.CFGERRUNCORIN(cfg_err_uncor_in)
   ,.CFGEXTFUNCTIONNUMBER(cfg_ext_function_number[7:0])
   ,.CFGEXTREADDATA(cfg_ext_read_data[31:0])
   ,.CFGEXTREADDATAVALID(cfg_ext_read_data_valid)
   ,.CFGEXTREADRECEIVED(cfg_ext_read_received)
   ,.CFGEXTREGISTERNUMBER(cfg_ext_register_number[9:0])
   ,.CFGEXTWRITEBYTEENABLE(cfg_ext_write_byte_enable[3:0])
   ,.CFGEXTWRITEDATA(cfg_ext_write_data[31:0])
   ,.CFGEXTWRITERECEIVED(cfg_ext_write_received)
   ,.CFGFCCPLD(cfg_fc_cpld[11:0])
   ,.CFGFCCPLH(cfg_fc_cplh[7:0])
   ,.CFGFCNPD(cfg_fc_npd[11:0])
   ,.CFGFCNPH(cfg_fc_nph[7:0])
   ,.CFGFCPD(cfg_fc_pd[11:0])
   ,.CFGFCPH(cfg_fc_ph[7:0])
   ,.CFGFCSEL(cfg_fc_sel[2:0])
   ,.CFGFLRDONE(cfg_flr_done[3:0])
   ,.CFGFLRINPROCESS(cfg_flr_in_process[3:0])
   ,.CFGFUNCTIONPOWERSTATE(cfg_function_power_state[11:0])
   ,.CFGFUNCTIONSTATUS(cfg_function_status[15:0])
   ,.CFGHOTRESETIN(cfg_hot_reset_in)
   ,.CFGHOTRESETOUT(cfg_hot_reset_out)
   ,.CFGINTERRUPTINT(cfg_interrupt_int[3:0])
   ,.CFGINTERRUPTMSIATTR(cfg_interrupt_msi_attr[2:0])
   ,.CFGINTERRUPTMSIDATA(cfg_interrupt_msi_data[31:0])
   ,.CFGINTERRUPTMSIENABLE(cfg_interrupt_msi_enable[3:0])
   ,.CFGINTERRUPTMSIFAIL(cfg_interrupt_msi_fail)
   ,.CFGINTERRUPTMSIFUNCTIONNUMBER(cfg_interrupt_msi_function_number[7:0])
   ,.CFGINTERRUPTMSIINT(cfg_interrupt_msi_int[31:0])
   ,.CFGINTERRUPTMSIMASKUPDATE(cfg_interrupt_msi_mask_update)
   ,.CFGINTERRUPTMSIMMENABLE(cfg_interrupt_msi_mmenable[11:0])
   ,.CFGINTERRUPTMSIPENDINGSTATUS(cfg_interrupt_msi_pending_status[31:0])
   ,.CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE(cfg_interrupt_msi_pending_status_data_enable)
   ,.CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM(cfg_interrupt_msi_pending_status_function_num[1:0])
   ,.CFGINTERRUPTMSISELECT(cfg_interrupt_msi_select[1:0])
   ,.CFGINTERRUPTMSISENT(cfg_interrupt_msi_sent)
   ,.CFGINTERRUPTMSITPHPRESENT(cfg_interrupt_msi_tph_present)
   ,.CFGINTERRUPTMSITPHSTTAG(cfg_interrupt_msi_tph_st_tag[7:0])
   ,.CFGINTERRUPTMSITPHTYPE(cfg_interrupt_msi_tph_type[1:0])
   ,.CFGINTERRUPTMSIXADDRESS(cfg_interrupt_msix_address[63:0])
   ,.CFGINTERRUPTMSIXDATA(cfg_interrupt_msix_data[31:0])
   ,.CFGINTERRUPTMSIXENABLE(cfg_interrupt_msix_enable[3:0])
   ,.CFGINTERRUPTMSIXINT(cfg_interrupt_msix_int)
   ,.CFGINTERRUPTMSIXMASK(cfg_interrupt_msix_mask[3:0])
   ,.CFGINTERRUPTMSIXVECPENDING(cfg_interrupt_msix_vec_pending[1:0])
   ,.CFGINTERRUPTMSIXVECPENDINGSTATUS(cfg_interrupt_msix_vec_pending_status)
   ,.CFGINTERRUPTPENDING(cfg_interrupt_pending[3:0])
   ,.CFGINTERRUPTSENT(cfg_interrupt_sent)
   ,.CFGLINKPOWERSTATE(cfg_link_power_state[1:0])
   ,.CFGLINKTRAININGENABLE(cfg_link_training_enable)
   ,.CFGLOCALERROROUT(cfg_local_error_out[4:0])
   ,.CFGLOCALERRORVALID(cfg_local_error_valid)
   ,.CFGLTRENABLE(cfg_ltr_enable)
   ,.CFGLTSSMSTATE(cfg_ltssm_state[5:0])
   ,.CFGMAXPAYLOAD(cfg_max_payload[1:0])
   ,.CFGMAXREADREQ(cfg_max_read_req[2:0])
   ,.CFGMGMTADDR(cfg_mgmt_addr[9:0])
   ,.CFGMGMTBYTEENABLE(cfg_mgmt_byte_enable[3:0])
   ,.CFGMGMTDEBUGACCESS(cfg_mgmt_debug_access)
   ,.CFGMGMTFUNCTIONNUMBER(cfg_mgmt_function_number[7:0])
   ,.CFGMGMTREAD(cfg_mgmt_read)
   ,.CFGMGMTREADDATA(cfg_mgmt_read_data[31:0])
   ,.CFGMGMTREADWRITEDONE(cfg_mgmt_read_write_done)
   ,.CFGMGMTWRITE(cfg_mgmt_write)
   ,.CFGMGMTWRITEDATA(cfg_mgmt_write_data[31:0])
   ,.CFGMSGRECEIVED(cfg_msg_received)
   ,.CFGMSGRECEIVEDDATA(cfg_msg_received_data[7:0])
   ,.CFGMSGRECEIVEDTYPE(cfg_msg_received_type[4:0])
   ,.CFGMSGTRANSMIT(cfg_msg_transmit)
   ,.CFGMSGTRANSMITDATA(cfg_msg_transmit_data[31:0])
   ,.CFGMSGTRANSMITDONE(cfg_msg_transmit_done)
   ,.CFGMSGTRANSMITTYPE(cfg_msg_transmit_type[2:0])
   ,.CFGMSIXRAMADDRESS(cfg_msix_ram_address[12:0])
   ,.CFGMSIXRAMREADDATA(cfg_msix_ram_read_data[35:0])
   ,.CFGMSIXRAMREADENABLE(cfg_msix_ram_read_enable)
   ,.CFGMSIXRAMWRITEBYTEENABLE(cfg_msix_ram_write_byte_enable[3:0])
   ,.CFGMSIXRAMWRITEDATA(cfg_msix_ram_write_data[35:0])
   ,.CFGNEGOTIATEDWIDTH(cfg_negotiated_width[2:0])
   ,.CFGOBFFENABLE(cfg_obff_enable[1:0])
   ,.CFGPHYLINKDOWN(cfg_phy_link_down_wire)
   ,.CFGPHYLINKSTATUS(cfg_phy_link_status[1:0])
   ,.CFGPLSTATUSCHANGE(cfg_pl_status_change)
   ,.CFGPMASPML1ENTRYREJECT(cfg_pm_aspm_l1_entry_reject)
   ,.CFGPMASPMTXL0SENTRYDISABLE(cfg_pm_aspm_tx_l0s_entry_disable)
   ,.CFGPOWERSTATECHANGEACK(cfg_power_state_change_ack)
   ,.CFGPOWERSTATECHANGEINTERRUPT(cfg_power_state_change_interrupt)
   ,.CFGRCBSTATUS(cfg_rcb_status[3:0])
   ,.CFGREQPMTRANSITIONL23READY(cfg_req_pm_transition_l23_ready)
   ,.CFGREVIDPF0(cfg_rev_id_pf0[7:0])
   ,.CFGREVIDPF1(cfg_rev_id_pf1[7:0])
   ,.CFGREVIDPF2(cfg_rev_id_pf2[7:0])
   ,.CFGREVIDPF3(cfg_rev_id_pf3[7:0])
   ,.CFGRXPMSTATE(cfg_rx_pm_state[1:0])
   ,.CFGSUBSYSIDPF0(cfg_subsys_id_pf0[15:0])
   ,.CFGSUBSYSIDPF1(cfg_subsys_id_pf1[15:0])
   ,.CFGSUBSYSIDPF2(cfg_subsys_id_pf2[15:0])
   ,.CFGSUBSYSIDPF3(cfg_subsys_id_pf3[15:0])
   ,.CFGSUBSYSVENDID(cfg_subsys_vend_id[15:0])
   ,.CFGTPHRAMADDRESS(cfg_tph_ram_address[11:0])
   ,.CFGTPHRAMREADDATA(cfg_tph_ram_read_data[35:0])
   ,.CFGTPHRAMREADENABLE(cfg_tph_ram_read_enable)
   ,.CFGTPHRAMWRITEBYTEENABLE(cfg_tph_ram_write_byte_enable[3:0])
   ,.CFGTPHRAMWRITEDATA(cfg_tph_ram_write_data[35:0])
   ,.CFGTPHREQUESTERENABLE(cfg_tph_requester_enable[3:0])
   ,.CFGTPHSTMODE(cfg_tph_st_mode[11:0])
   ,.CFGTXPMSTATE(cfg_tx_pm_state[1:0])
   ,.CFGVENDID(cfg_vend_id[15:0])
   ,.CFGVFFLRDONE(cfg_vf_flr_done)
   ,.CFGVFFLRFUNCNUM(cfg_vf_flr_func_num[7:0])
   ,.CONFMCAPDESIGNSWITCH(conf_mcap_design_switch)
   ,.CONFMCAPEOS(conf_mcap_eos)
   ,.CONFMCAPINUSEBYPCIE(conf_mcap_in_use_by_pcie)
   ,.CONFMCAPREQUESTBYCONF(conf_mcap_request_by_conf)
   ,.CONFREQDATA(conf_req_data[31:0])
   ,.CONFREQREADY(conf_req_ready)
   ,.CONFREQREGNUM(conf_req_reg_num[3:0])
   ,.CONFREQTYPE(conf_req_type[1:0])
   ,.CONFREQVALID(conf_req_valid)
   ,.CONFRESPRDATA(conf_resp_rdata[31:0])
   ,.CONFRESPVALID(conf_resp_valid)
   ,.CORECLK(core_clk)
   ,.CORECLKMIREPLAYRAM0(core_clk)
   ,.CORECLKMIREPLAYRAM1(core_clk)
   ,.CORECLKMIRXCOMPLETIONRAM0(core_clk)
   ,.CORECLKMIRXCOMPLETIONRAM1(core_clk)
   ,.CORECLKMIRXPOSTEDREQUESTRAM0(core_clk)
   ,.CORECLKMIRXPOSTEDREQUESTRAM1(core_clk)
   ,.DBGCTRL0OUT( )
   ,.DBGCTRL1OUT( )
   ,.DBGDATA0OUT( )
   ,.DBGDATA1OUT( )
   ,.DBGSEL0(6'd0)
   ,.DBGSEL1(6'd0)
   ,.DRPADDR(drp_addr[9:0])
   ,.DRPCLK(drp_clk)
   ,.DRPDI(drp_di[15:0])
   ,.DRPDO(drp_do[15:0])
   ,.DRPEN(drp_en)
   ,.DRPRDY(drp_rdy)
   ,.DRPWE(drp_we)
   ,.MAXISCQTDATA(m_axis_cq_tdata_int[255:0])
   ,.MAXISCQTKEEP(m_axis_cq_tkeep_int[7:0])
   ,.MAXISCQTLAST(m_axis_cq_tlast_int)
   ,.MAXISCQTREADY(m_axis_cq_tready_int[21:0])
   ,.MAXISCQTUSER(m_axis_cq_tuser_int[87:0])
   ,.MAXISCQTVALID(m_axis_cq_tvalid_int)
   ,.MAXISRCTDATA(m_axis_rc_tdata_int[255:0])
   ,.MAXISRCTKEEP(m_axis_rc_tkeep_int[7:0])
   ,.MAXISRCTLAST(m_axis_rc_tlast_int)
   ,.MAXISRCTREADY(m_axis_rc_tready_int[21:0])
   ,.MAXISRCTUSER(m_axis_rc_tuser_int[74:0])
   ,.MAXISRCTVALID(m_axis_rc_tvalid_int)
   ,.MCAPCLK(mcap_clk)
   ,.MGMTRESETN(mgmt_reset_n)
   ,.MGMTSTICKYRESETN(mgmt_sticky_reset_n)
   ,.MIREPLAYRAMADDRESS0(mi_replay_ram_address0[8:0])
   ,.MIREPLAYRAMADDRESS1(mi_replay_ram_address1[8:0])
   ,.MIREPLAYRAMERRCOR(mi_replay_ram_err_cor[5:0])
   ,.MIREPLAYRAMERRUNCOR(mi_replay_ram_err_uncor[5:0])
   ,.MIREPLAYRAMREADDATA0(mi_replay_ram_read_data0[127:0])
   ,.MIREPLAYRAMREADDATA1(mi_replay_ram_read_data1[127:0])
   ,.MIREPLAYRAMREADENABLE0(mi_replay_ram_read_enable0)
   ,.MIREPLAYRAMREADENABLE1(mi_replay_ram_read_enable1)
   ,.MIREPLAYRAMWRITEDATA0(mi_replay_ram_write_data0[127:0])
   ,.MIREPLAYRAMWRITEDATA1(mi_replay_ram_write_data1[127:0])
   ,.MIREPLAYRAMWRITEENABLE0(mi_replay_ram_write_enable0)
   ,.MIREPLAYRAMWRITEENABLE1(mi_replay_ram_write_enable1)
   ,.MIRXCOMPLETIONRAMERRCOR(mi_rx_completion_ram_err_cor[11:0])
   ,.MIRXCOMPLETIONRAMERRUNCOR(mi_rx_completion_ram_err_uncor[11:0])
   ,.MIRXCOMPLETIONRAMREADADDRESS0(mi_rx_completion_ram_read_address0[8:0])
   ,.MIRXCOMPLETIONRAMREADADDRESS1(mi_rx_completion_ram_read_address1[8:0])
   ,.MIRXCOMPLETIONRAMREADDATA0(mi_rx_completion_ram_read_data0[143:0])
   ,.MIRXCOMPLETIONRAMREADDATA1(mi_rx_completion_ram_read_data1[143:0])
   ,.MIRXCOMPLETIONRAMREADENABLE0(mi_rx_completion_ram_read_enable0[1:0])
   ,.MIRXCOMPLETIONRAMREADENABLE1(mi_rx_completion_ram_read_enable1[1:0])
   ,.MIRXCOMPLETIONRAMWRITEADDRESS0(mi_rx_completion_ram_write_address0[8:0])
   ,.MIRXCOMPLETIONRAMWRITEADDRESS1(mi_rx_completion_ram_write_address1[8:0])
   ,.MIRXCOMPLETIONRAMWRITEDATA0(mi_rx_completion_ram_write_data0[143:0])
   ,.MIRXCOMPLETIONRAMWRITEDATA1(mi_rx_completion_ram_write_data1[143:0])
   ,.MIRXCOMPLETIONRAMWRITEENABLE0(mi_rx_completion_ram_write_enable0[1:0])
   ,.MIRXCOMPLETIONRAMWRITEENABLE1(mi_rx_completion_ram_write_enable1[1:0])
   ,.MIRXPOSTEDREQUESTRAMERRCOR(mi_rx_posted_request_ram_err_cor[5:0])
   ,.MIRXPOSTEDREQUESTRAMERRUNCOR(mi_rx_posted_request_ram_err_uncor[5:0])
   ,.MIRXPOSTEDREQUESTRAMREADADDRESS0(mi_rx_posted_request_ram_read_address0[8:0])
   ,.MIRXPOSTEDREQUESTRAMREADADDRESS1(mi_rx_posted_request_ram_read_address1[8:0])
   ,.MIRXPOSTEDREQUESTRAMREADDATA0(mi_rx_posted_request_ram_read_data0[143:0])
   ,.MIRXPOSTEDREQUESTRAMREADDATA1(mi_rx_posted_request_ram_read_data1[143:0])
   ,.MIRXPOSTEDREQUESTRAMREADENABLE0(mi_rx_posted_request_ram_read_enable0)
   ,.MIRXPOSTEDREQUESTRAMREADENABLE1(mi_rx_posted_request_ram_read_enable1)
   ,.MIRXPOSTEDREQUESTRAMWRITEADDRESS0(mi_rx_posted_request_ram_write_address0[8:0])
   ,.MIRXPOSTEDREQUESTRAMWRITEADDRESS1(mi_rx_posted_request_ram_write_address1[8:0])
   ,.MIRXPOSTEDREQUESTRAMWRITEDATA0(mi_rx_posted_request_ram_write_data0[143:0])
   ,.MIRXPOSTEDREQUESTRAMWRITEDATA1(mi_rx_posted_request_ram_write_data1[143:0])
   ,.MIRXPOSTEDREQUESTRAMWRITEENABLE0(mi_rx_posted_request_ram_write_enable0)
   ,.MIRXPOSTEDREQUESTRAMWRITEENABLE1(mi_rx_posted_request_ram_write_enable1)
   ,.PCIECOMPLDELIVERED(pcie_compl_delivered[1:0])
   ,.PCIECOMPLDELIVEREDTAG0(pcie_compl_delivered_tag0[7:0])
   ,.PCIECOMPLDELIVEREDTAG1(pcie_compl_delivered_tag1[7:0])
   ,.PCIECQNPREQ(pcie_cq_np_req[1:0])
   ,.PCIECQNPREQCOUNT(pcie_cq_np_req_count_int[5:0])
   ,.PCIECQNPUSERCREDITRCVD(pcie_cq_np_user_credit_rcvd)
   ,.PCIECQPIPELINEEMPTY(pcie_cq_pipeline_empty)
   ,.PCIEPERST0B(pcie_perst0_b)
   ,.PCIEPERST1B(pcie_perst1_b)
   ,.MCAPPERST0B(mcap_rst_b)
   ,.MCAPPERST1B(mcap_rst_b)
   ,.PCIEPOSTEDREQDELIVERED(pcie_posted_req_delivered)
   ,.PCIERQSEQNUM0(pcie_rq_seq_num0_cc[5:0])
   ,.PCIERQSEQNUM1(pcie_rq_seq_num1[5:0])
   ,.PCIERQSEQNUMVLD0(pcie_rq_seq_num_vld0_cc)
   ,.PCIERQSEQNUMVLD1(pcie_rq_seq_num_vld1)
   ,.PCIERQTAG0(pcie_rq_tag0[7:0])
   ,.PCIERQTAG1(pcie_rq_tag1[7:0])
   ,.PCIERQTAGAV(pcie_rq_tag_av[3:0])
   ,.PCIERQTAGVLD0(pcie_rq_tag_vld0)
   ,.PCIERQTAGVLD1(pcie_rq_tag_vld1)
   ,.PCIETFCNPDAV(pcie_tfc_npd_av[3:0])
   ,.PCIETFCNPHAV(pcie_tfc_nph_av[3:0])
   ,.PIPECLKEN(1'b1)
   ,.PIPECLK(pipe_clk_to_e4)
   ,.PIPEEQFS(pipe_eq_fs[5:0])
   ,.PIPEEQLF(pipe_eq_lf[5:0])
   ,.PIPERESETN(pipe_reset_n)
   ,.PIPERX00CHARISK(pipe_rx00_char_is_k[1:0])
   ,.PIPERX00DATA(pipe_rx00_data[31:0])
   ,.PIPERX00DATAVALID(pipe_rx00_data_valid)
   ,.PIPERX00ELECIDLE(pipe_rx00_elec_idle)
   ,.PIPERX00EQCONTROL(pipe_rx00_eq_control[1:0])
   ,.PIPERX00EQDONE(pipe_rx00_eq_done)
   ,.PIPERX00EQLPADAPTDONE(pipe_rx00_eq_lp_adapt_done)
   ,.PIPERX00EQLPLFFSSEL(pipe_rx00_eq_lp_lf_fs_sel)
   ,.PIPERX00EQLPNEWTXCOEFFORPRESET(pipe_rx00_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX00PHYSTATUS(pipe_rx00_phy_status)
   ,.PIPERX00POLARITY(pipe_rx00_polarity)
   ,.PIPERX00STARTBLOCK(pipe_rx00_start_block[1:0])
   ,.PIPERX00STATUS(pipe_rx00_status[2:0])
   ,.PIPERX00SYNCHEADER(pipe_rx00_sync_header[1:0])
   ,.PIPERX00VALID(pipe_rx00_valid)
   ,.PIPERX01CHARISK(pipe_rx01_char_is_k[1:0])
   ,.PIPERX01DATA(pipe_rx01_data[31:0])
   ,.PIPERX01DATAVALID(pipe_rx01_data_valid)
   ,.PIPERX01ELECIDLE(pipe_rx01_elec_idle)
   ,.PIPERX01EQCONTROL(pipe_rx01_eq_control[1:0])
   ,.PIPERX01EQDONE(pipe_rx01_eq_done)
   ,.PIPERX01EQLPADAPTDONE(pipe_rx01_eq_lp_adapt_done)
   ,.PIPERX01EQLPLFFSSEL(pipe_rx01_eq_lp_lf_fs_sel)
   ,.PIPERX01EQLPNEWTXCOEFFORPRESET(pipe_rx01_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX01PHYSTATUS(pipe_rx01_phy_status)
   ,.PIPERX01POLARITY(pipe_rx01_polarity)
   ,.PIPERX01STARTBLOCK(pipe_rx01_start_block[1:0])
   ,.PIPERX01STATUS(pipe_rx01_status[2:0])
   ,.PIPERX01SYNCHEADER(pipe_rx01_sync_header[1:0])
   ,.PIPERX01VALID(pipe_rx01_valid)
   ,.PIPERX02CHARISK(pipe_rx02_char_is_k[1:0])
   ,.PIPERX02DATA(pipe_rx02_data[31:0])
   ,.PIPERX02DATAVALID(pipe_rx02_data_valid)
   ,.PIPERX02ELECIDLE(pipe_rx02_elec_idle)
   ,.PIPERX02EQCONTROL(pipe_rx02_eq_control[1:0])
   ,.PIPERX02EQDONE(pipe_rx02_eq_done)
   ,.PIPERX02EQLPADAPTDONE(pipe_rx02_eq_lp_adapt_done)
   ,.PIPERX02EQLPLFFSSEL(pipe_rx02_eq_lp_lf_fs_sel)
   ,.PIPERX02EQLPNEWTXCOEFFORPRESET(pipe_rx02_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX02PHYSTATUS(pipe_rx02_phy_status)
   ,.PIPERX02POLARITY(pipe_rx02_polarity)
   ,.PIPERX02STARTBLOCK(pipe_rx02_start_block[1:0])
   ,.PIPERX02STATUS(pipe_rx02_status[2:0])
   ,.PIPERX02SYNCHEADER(pipe_rx02_sync_header[1:0])
   ,.PIPERX02VALID(pipe_rx02_valid)
   ,.PIPERX03CHARISK(pipe_rx03_char_is_k[1:0])
   ,.PIPERX03DATA(pipe_rx03_data[31:0])
   ,.PIPERX03DATAVALID(pipe_rx03_data_valid)
   ,.PIPERX03ELECIDLE(pipe_rx03_elec_idle)
   ,.PIPERX03EQCONTROL(pipe_rx03_eq_control[1:0])
   ,.PIPERX03EQDONE(pipe_rx03_eq_done)
   ,.PIPERX03EQLPADAPTDONE(pipe_rx03_eq_lp_adapt_done)
   ,.PIPERX03EQLPLFFSSEL(pipe_rx03_eq_lp_lf_fs_sel)
   ,.PIPERX03EQLPNEWTXCOEFFORPRESET(pipe_rx03_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX03PHYSTATUS(pipe_rx03_phy_status)
   ,.PIPERX03POLARITY(pipe_rx03_polarity)
   ,.PIPERX03STARTBLOCK(pipe_rx03_start_block[1:0])
   ,.PIPERX03STATUS(pipe_rx03_status[2:0])
   ,.PIPERX03SYNCHEADER(pipe_rx03_sync_header[1:0])
   ,.PIPERX03VALID(pipe_rx03_valid)
   ,.PIPERX04CHARISK(pipe_rx04_char_is_k[1:0])
   ,.PIPERX04DATA(pipe_rx04_data[31:0])
   ,.PIPERX04DATAVALID(pipe_rx04_data_valid)
   ,.PIPERX04ELECIDLE(pipe_rx04_elec_idle)
   ,.PIPERX04EQCONTROL(pipe_rx04_eq_control[1:0])
   ,.PIPERX04EQDONE(pipe_rx04_eq_done)
   ,.PIPERX04EQLPADAPTDONE(pipe_rx04_eq_lp_adapt_done)
   ,.PIPERX04EQLPLFFSSEL(pipe_rx04_eq_lp_lf_fs_sel)
   ,.PIPERX04EQLPNEWTXCOEFFORPRESET(pipe_rx04_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX04PHYSTATUS(pipe_rx04_phy_status)
   ,.PIPERX04POLARITY(pipe_rx04_polarity)
   ,.PIPERX04STARTBLOCK(pipe_rx04_start_block[1:0])
   ,.PIPERX04STATUS(pipe_rx04_status[2:0])
   ,.PIPERX04SYNCHEADER(pipe_rx04_sync_header[1:0])
   ,.PIPERX04VALID(pipe_rx04_valid)
   ,.PIPERX05CHARISK(pipe_rx05_char_is_k[1:0])
   ,.PIPERX05DATA(pipe_rx05_data[31:0])
   ,.PIPERX05DATAVALID(pipe_rx05_data_valid)
   ,.PIPERX05ELECIDLE(pipe_rx05_elec_idle)
   ,.PIPERX05EQCONTROL(pipe_rx05_eq_control[1:0])
   ,.PIPERX05EQDONE(pipe_rx05_eq_done)
   ,.PIPERX05EQLPADAPTDONE(pipe_rx05_eq_lp_adapt_done)
   ,.PIPERX05EQLPLFFSSEL(pipe_rx05_eq_lp_lf_fs_sel)
   ,.PIPERX05EQLPNEWTXCOEFFORPRESET(pipe_rx05_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX05PHYSTATUS(pipe_rx05_phy_status)
   ,.PIPERX05POLARITY(pipe_rx05_polarity)
   ,.PIPERX05STARTBLOCK(pipe_rx05_start_block[1:0])
   ,.PIPERX05STATUS(pipe_rx05_status[2:0])
   ,.PIPERX05SYNCHEADER(pipe_rx05_sync_header[1:0])
   ,.PIPERX05VALID(pipe_rx05_valid)
   ,.PIPERX06CHARISK(pipe_rx06_char_is_k[1:0])
   ,.PIPERX06DATA(pipe_rx06_data[31:0])
   ,.PIPERX06DATAVALID(pipe_rx06_data_valid)
   ,.PIPERX06ELECIDLE(pipe_rx06_elec_idle)
   ,.PIPERX06EQCONTROL(pipe_rx06_eq_control[1:0])
   ,.PIPERX06EQDONE(pipe_rx06_eq_done)
   ,.PIPERX06EQLPADAPTDONE(pipe_rx06_eq_lp_adapt_done)
   ,.PIPERX06EQLPLFFSSEL(pipe_rx06_eq_lp_lf_fs_sel)
   ,.PIPERX06EQLPNEWTXCOEFFORPRESET(pipe_rx06_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX06PHYSTATUS(pipe_rx06_phy_status)
   ,.PIPERX06POLARITY(pipe_rx06_polarity)
   ,.PIPERX06STARTBLOCK(pipe_rx06_start_block[1:0])
   ,.PIPERX06STATUS(pipe_rx06_status[2:0])
   ,.PIPERX06SYNCHEADER(pipe_rx06_sync_header[1:0])
   ,.PIPERX06VALID(pipe_rx06_valid)
   ,.PIPERX07CHARISK(pipe_rx07_char_is_k[1:0])
   ,.PIPERX07DATA(pipe_rx07_data[31:0])
   ,.PIPERX07DATAVALID(pipe_rx07_data_valid)
   ,.PIPERX07ELECIDLE(pipe_rx07_elec_idle)
   ,.PIPERX07EQCONTROL(pipe_rx07_eq_control[1:0])
   ,.PIPERX07EQDONE(pipe_rx07_eq_done)
   ,.PIPERX07EQLPADAPTDONE(pipe_rx07_eq_lp_adapt_done)
   ,.PIPERX07EQLPLFFSSEL(pipe_rx07_eq_lp_lf_fs_sel)
   ,.PIPERX07EQLPNEWTXCOEFFORPRESET(pipe_rx07_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX07PHYSTATUS(pipe_rx07_phy_status)
   ,.PIPERX07POLARITY(pipe_rx07_polarity)
   ,.PIPERX07STARTBLOCK(pipe_rx07_start_block[1:0])
   ,.PIPERX07STATUS(pipe_rx07_status[2:0])
   ,.PIPERX07SYNCHEADER(pipe_rx07_sync_header[1:0])
   ,.PIPERX07VALID(pipe_rx07_valid)
   ,.PIPERX08CHARISK(pipe_rx08_char_is_k[1:0])
   ,.PIPERX08DATA(pipe_rx08_data[31:0])
   ,.PIPERX08DATAVALID(pipe_rx08_data_valid)
   ,.PIPERX08ELECIDLE(pipe_rx08_elec_idle)
   ,.PIPERX08EQCONTROL(pipe_rx08_eq_control[1:0])
   ,.PIPERX08EQDONE(pipe_rx08_eq_done)
   ,.PIPERX08EQLPADAPTDONE(pipe_rx08_eq_lp_adapt_done)
   ,.PIPERX08EQLPLFFSSEL(pipe_rx08_eq_lp_lf_fs_sel)
   ,.PIPERX08EQLPNEWTXCOEFFORPRESET(pipe_rx08_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX08PHYSTATUS(pipe_rx08_phy_status)
   ,.PIPERX08POLARITY(pipe_rx08_polarity)
   ,.PIPERX08STARTBLOCK(pipe_rx08_start_block[1:0])
   ,.PIPERX08STATUS(pipe_rx08_status[2:0])
   ,.PIPERX08SYNCHEADER(pipe_rx08_sync_header[1:0])
   ,.PIPERX08VALID(pipe_rx08_valid)
   ,.PIPERX09CHARISK(pipe_rx09_char_is_k[1:0])
   ,.PIPERX09DATA(pipe_rx09_data[31:0])
   ,.PIPERX09DATAVALID(pipe_rx09_data_valid)
   ,.PIPERX09ELECIDLE(pipe_rx09_elec_idle)
   ,.PIPERX09EQCONTROL(pipe_rx09_eq_control[1:0])
   ,.PIPERX09EQDONE(pipe_rx09_eq_done)
   ,.PIPERX09EQLPADAPTDONE(pipe_rx09_eq_lp_adapt_done)
   ,.PIPERX09EQLPLFFSSEL(pipe_rx09_eq_lp_lf_fs_sel)
   ,.PIPERX09EQLPNEWTXCOEFFORPRESET(pipe_rx09_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX09PHYSTATUS(pipe_rx09_phy_status)
   ,.PIPERX09POLARITY(pipe_rx09_polarity)
   ,.PIPERX09STARTBLOCK(pipe_rx09_start_block[1:0])
   ,.PIPERX09STATUS(pipe_rx09_status[2:0])
   ,.PIPERX09SYNCHEADER(pipe_rx09_sync_header[1:0])
   ,.PIPERX09VALID(pipe_rx09_valid)
   ,.PIPERX10CHARISK(pipe_rx10_char_is_k[1:0])
   ,.PIPERX10DATA(pipe_rx10_data[31:0])
   ,.PIPERX10DATAVALID(pipe_rx10_data_valid)
   ,.PIPERX10ELECIDLE(pipe_rx10_elec_idle)
   ,.PIPERX10EQCONTROL(pipe_rx10_eq_control[1:0])
   ,.PIPERX10EQDONE(pipe_rx10_eq_done)
   ,.PIPERX10EQLPADAPTDONE(pipe_rx10_eq_lp_adapt_done)
   ,.PIPERX10EQLPLFFSSEL(pipe_rx10_eq_lp_lf_fs_sel)
   ,.PIPERX10EQLPNEWTXCOEFFORPRESET(pipe_rx10_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX10PHYSTATUS(pipe_rx10_phy_status)
   ,.PIPERX10POLARITY(pipe_rx10_polarity)
   ,.PIPERX10STARTBLOCK(pipe_rx10_start_block[1:0])
   ,.PIPERX10STATUS(pipe_rx10_status[2:0])
   ,.PIPERX10SYNCHEADER(pipe_rx10_sync_header[1:0])
   ,.PIPERX10VALID(pipe_rx10_valid)
   ,.PIPERX11CHARISK(pipe_rx11_char_is_k[1:0])
   ,.PIPERX11DATA(pipe_rx11_data[31:0])
   ,.PIPERX11DATAVALID(pipe_rx11_data_valid)
   ,.PIPERX11ELECIDLE(pipe_rx11_elec_idle)
   ,.PIPERX11EQCONTROL(pipe_rx11_eq_control[1:0])
   ,.PIPERX11EQDONE(pipe_rx11_eq_done)
   ,.PIPERX11EQLPADAPTDONE(pipe_rx11_eq_lp_adapt_done)
   ,.PIPERX11EQLPLFFSSEL(pipe_rx11_eq_lp_lf_fs_sel)
   ,.PIPERX11EQLPNEWTXCOEFFORPRESET(pipe_rx11_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX11PHYSTATUS(pipe_rx11_phy_status)
   ,.PIPERX11POLARITY(pipe_rx11_polarity)
   ,.PIPERX11STARTBLOCK(pipe_rx11_start_block[1:0])
   ,.PIPERX11STATUS(pipe_rx11_status[2:0])
   ,.PIPERX11SYNCHEADER(pipe_rx11_sync_header[1:0])
   ,.PIPERX11VALID(pipe_rx11_valid)
   ,.PIPERX12CHARISK(pipe_rx12_char_is_k[1:0])
   ,.PIPERX12DATA(pipe_rx12_data[31:0])
   ,.PIPERX12DATAVALID(pipe_rx12_data_valid)
   ,.PIPERX12ELECIDLE(pipe_rx12_elec_idle)
   ,.PIPERX12EQCONTROL(pipe_rx12_eq_control[1:0])
   ,.PIPERX12EQDONE(pipe_rx12_eq_done)
   ,.PIPERX12EQLPADAPTDONE(pipe_rx12_eq_lp_adapt_done)
   ,.PIPERX12EQLPLFFSSEL(pipe_rx12_eq_lp_lf_fs_sel)
   ,.PIPERX12EQLPNEWTXCOEFFORPRESET(pipe_rx12_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX12PHYSTATUS(pipe_rx12_phy_status)
   ,.PIPERX12POLARITY(pipe_rx12_polarity)
   ,.PIPERX12STARTBLOCK(pipe_rx12_start_block[1:0])
   ,.PIPERX12STATUS(pipe_rx12_status[2:0])
   ,.PIPERX12SYNCHEADER(pipe_rx12_sync_header[1:0])
   ,.PIPERX12VALID(pipe_rx12_valid)
   ,.PIPERX13CHARISK(pipe_rx13_char_is_k[1:0])
   ,.PIPERX13DATA(pipe_rx13_data[31:0])
   ,.PIPERX13DATAVALID(pipe_rx13_data_valid)
   ,.PIPERX13ELECIDLE(pipe_rx13_elec_idle)
   ,.PIPERX13EQCONTROL(pipe_rx13_eq_control[1:0])
   ,.PIPERX13EQDONE(pipe_rx13_eq_done)
   ,.PIPERX13EQLPADAPTDONE(pipe_rx13_eq_lp_adapt_done)
   ,.PIPERX13EQLPLFFSSEL(pipe_rx13_eq_lp_lf_fs_sel)
   ,.PIPERX13EQLPNEWTXCOEFFORPRESET(pipe_rx13_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX13PHYSTATUS(pipe_rx13_phy_status)
   ,.PIPERX13POLARITY(pipe_rx13_polarity)
   ,.PIPERX13STARTBLOCK(pipe_rx13_start_block[1:0])
   ,.PIPERX13STATUS(pipe_rx13_status[2:0])
   ,.PIPERX13SYNCHEADER(pipe_rx13_sync_header[1:0])
   ,.PIPERX13VALID(pipe_rx13_valid)
   ,.PIPERX14CHARISK(pipe_rx14_char_is_k[1:0])
   ,.PIPERX14DATA(pipe_rx14_data[31:0])
   ,.PIPERX14DATAVALID(pipe_rx14_data_valid)
   ,.PIPERX14ELECIDLE(pipe_rx14_elec_idle)
   ,.PIPERX14EQCONTROL(pipe_rx14_eq_control[1:0])
   ,.PIPERX14EQDONE(pipe_rx14_eq_done)
   ,.PIPERX14EQLPADAPTDONE(pipe_rx14_eq_lp_adapt_done)
   ,.PIPERX14EQLPLFFSSEL(pipe_rx14_eq_lp_lf_fs_sel)
   ,.PIPERX14EQLPNEWTXCOEFFORPRESET(pipe_rx14_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX14PHYSTATUS(pipe_rx14_phy_status)
   ,.PIPERX14POLARITY(pipe_rx14_polarity)
   ,.PIPERX14STARTBLOCK(pipe_rx14_start_block[1:0])
   ,.PIPERX14STATUS(pipe_rx14_status[2:0])
   ,.PIPERX14SYNCHEADER(pipe_rx14_sync_header[1:0])
   ,.PIPERX14VALID(pipe_rx14_valid)
   ,.PIPERX15CHARISK(pipe_rx15_char_is_k[1:0])
   ,.PIPERX15DATA(pipe_rx15_data[31:0])
   ,.PIPERX15DATAVALID(pipe_rx15_data_valid)
   ,.PIPERX15ELECIDLE(pipe_rx15_elec_idle)
   ,.PIPERX15EQCONTROL(pipe_rx15_eq_control[1:0])
   ,.PIPERX15EQDONE(pipe_rx15_eq_done)
   ,.PIPERX15EQLPADAPTDONE(pipe_rx15_eq_lp_adapt_done)
   ,.PIPERX15EQLPLFFSSEL(pipe_rx15_eq_lp_lf_fs_sel)
   ,.PIPERX15EQLPNEWTXCOEFFORPRESET(pipe_rx15_eq_lp_new_tx_coeff_or_preset[17:0])
   ,.PIPERX15PHYSTATUS(pipe_rx15_phy_status)
   ,.PIPERX15POLARITY(pipe_rx15_polarity)
   ,.PIPERX15STARTBLOCK(pipe_rx15_start_block[1:0])
   ,.PIPERX15STATUS(pipe_rx15_status[2:0])
   ,.PIPERX15SYNCHEADER(pipe_rx15_sync_header[1:0])
   ,.PIPERX15VALID(pipe_rx15_valid)
   ,.PIPERXEQLPLFFS(pipe_rx_eq_lp_lf_fs[5:0])
   ,.PIPERXEQLPTXPRESET(pipe_rx_eq_lp_tx_preset[3:0])
   ,.PIPETX00CHARISK(pipe_tx00_char_is_k[1:0])
   ,.PIPETX00COMPLIANCE(pipe_tx00_compliance)
   ,.PIPETX00DATA(pipe_tx00_data_out[31:0])
   ,.PIPETX00DATAVALID(pipe_tx00_data_valid)
   ,.PIPETX00ELECIDLE(pipe_tx00_elec_idle)
   ,.PIPETX00EQCOEFF(pipe_tx00_eq_coeff[17:0])
   ,.PIPETX00EQCONTROL(pipe_tx00_eq_control[1:0])
   ,.PIPETX00EQDEEMPH(pipe_tx00_eq_deemph[5:0])
   ,.PIPETX00EQDONE(pipe_tx00_eq_done)
   ,.PIPETX00POWERDOWN(pipe_tx00_powerdown[1:0])
   ,.PIPETX00STARTBLOCK(pipe_tx00_start_block)
   ,.PIPETX00SYNCHEADER(pipe_tx00_sync_header[1:0])
   ,.PIPETX01CHARISK(pipe_tx01_char_is_k[1:0])
   ,.PIPETX01COMPLIANCE(pipe_tx01_compliance)
   ,.PIPETX01DATA(pipe_tx01_data_out[31:0])
   ,.PIPETX01DATAVALID(pipe_tx01_data_valid)
   ,.PIPETX01ELECIDLE(pipe_tx01_elec_idle)
   ,.PIPETX01EQCOEFF(pipe_tx01_eq_coeff[17:0])
   ,.PIPETX01EQCONTROL(pipe_tx01_eq_control[1:0])
   ,.PIPETX01EQDEEMPH(pipe_tx01_eq_deemph[5:0])
   ,.PIPETX01EQDONE(pipe_tx01_eq_done)
   ,.PIPETX01POWERDOWN(pipe_tx01_powerdown[1:0])
   ,.PIPETX01STARTBLOCK(pipe_tx01_start_block)
   ,.PIPETX01SYNCHEADER(pipe_tx01_sync_header[1:0])
   ,.PIPETX02CHARISK(pipe_tx02_char_is_k[1:0])
   ,.PIPETX02COMPLIANCE(pipe_tx02_compliance)
   ,.PIPETX02DATA(pipe_tx02_data_out[31:0])
   ,.PIPETX02DATAVALID(pipe_tx02_data_valid)
   ,.PIPETX02ELECIDLE(pipe_tx02_elec_idle)
   ,.PIPETX02EQCOEFF(pipe_tx02_eq_coeff[17:0])
   ,.PIPETX02EQCONTROL(pipe_tx02_eq_control[1:0])
   ,.PIPETX02EQDEEMPH(pipe_tx02_eq_deemph[5:0])
   ,.PIPETX02EQDONE(pipe_tx02_eq_done)
   ,.PIPETX02POWERDOWN(pipe_tx02_powerdown[1:0])
   ,.PIPETX02STARTBLOCK(pipe_tx02_start_block)
   ,.PIPETX02SYNCHEADER(pipe_tx02_sync_header[1:0])
   ,.PIPETX03CHARISK(pipe_tx03_char_is_k[1:0])
   ,.PIPETX03COMPLIANCE(pipe_tx03_compliance)
   ,.PIPETX03DATA(pipe_tx03_data_out[31:0])
   ,.PIPETX03DATAVALID(pipe_tx03_data_valid)
   ,.PIPETX03ELECIDLE(pipe_tx03_elec_idle)
   ,.PIPETX03EQCOEFF(pipe_tx03_eq_coeff[17:0])
   ,.PIPETX03EQCONTROL(pipe_tx03_eq_control[1:0])
   ,.PIPETX03EQDEEMPH(pipe_tx03_eq_deemph[5:0])
   ,.PIPETX03EQDONE(pipe_tx03_eq_done)
   ,.PIPETX03POWERDOWN(pipe_tx03_powerdown[1:0])
   ,.PIPETX03STARTBLOCK(pipe_tx03_start_block)
   ,.PIPETX03SYNCHEADER(pipe_tx03_sync_header[1:0])
   ,.PIPETX04CHARISK(pipe_tx04_char_is_k[1:0])
   ,.PIPETX04COMPLIANCE(pipe_tx04_compliance)
   ,.PIPETX04DATA(pipe_tx04_data_out[31:0])
   ,.PIPETX04DATAVALID(pipe_tx04_data_valid)
   ,.PIPETX04ELECIDLE(pipe_tx04_elec_idle)
   ,.PIPETX04EQCOEFF(pipe_tx04_eq_coeff[17:0])
   ,.PIPETX04EQCONTROL(pipe_tx04_eq_control[1:0])
   ,.PIPETX04EQDEEMPH(pipe_tx04_eq_deemph[5:0])
   ,.PIPETX04EQDONE(pipe_tx04_eq_done)
   ,.PIPETX04POWERDOWN(pipe_tx04_powerdown[1:0])
   ,.PIPETX04STARTBLOCK(pipe_tx04_start_block)
   ,.PIPETX04SYNCHEADER(pipe_tx04_sync_header[1:0])
   ,.PIPETX05CHARISK(pipe_tx05_char_is_k[1:0])
   ,.PIPETX05COMPLIANCE(pipe_tx05_compliance)
   ,.PIPETX05DATA(pipe_tx05_data_out[31:0])
   ,.PIPETX05DATAVALID(pipe_tx05_data_valid)
   ,.PIPETX05ELECIDLE(pipe_tx05_elec_idle)
   ,.PIPETX05EQCOEFF(pipe_tx05_eq_coeff[17:0])
   ,.PIPETX05EQCONTROL(pipe_tx05_eq_control[1:0])
   ,.PIPETX05EQDEEMPH(pipe_tx05_eq_deemph[5:0])
   ,.PIPETX05EQDONE(pipe_tx05_eq_done)
   ,.PIPETX05POWERDOWN(pipe_tx05_powerdown[1:0])
   ,.PIPETX05STARTBLOCK(pipe_tx05_start_block)
   ,.PIPETX05SYNCHEADER(pipe_tx05_sync_header[1:0])
   ,.PIPETX06CHARISK(pipe_tx06_char_is_k[1:0])
   ,.PIPETX06COMPLIANCE(pipe_tx06_compliance)
   ,.PIPETX06DATA(pipe_tx06_data_out[31:0])
   ,.PIPETX06DATAVALID(pipe_tx06_data_valid)
   ,.PIPETX06ELECIDLE(pipe_tx06_elec_idle)
   ,.PIPETX06EQCOEFF(pipe_tx06_eq_coeff[17:0])
   ,.PIPETX06EQCONTROL(pipe_tx06_eq_control[1:0])
   ,.PIPETX06EQDEEMPH(pipe_tx06_eq_deemph[5:0])
   ,.PIPETX06EQDONE(pipe_tx06_eq_done)
   ,.PIPETX06POWERDOWN(pipe_tx06_powerdown[1:0])
   ,.PIPETX06STARTBLOCK(pipe_tx06_start_block)
   ,.PIPETX06SYNCHEADER(pipe_tx06_sync_header[1:0])
   ,.PIPETX07CHARISK(pipe_tx07_char_is_k[1:0])
   ,.PIPETX07COMPLIANCE(pipe_tx07_compliance)
   ,.PIPETX07DATA(pipe_tx07_data_out[31:0])
   ,.PIPETX07DATAVALID(pipe_tx07_data_valid)
   ,.PIPETX07ELECIDLE(pipe_tx07_elec_idle)
   ,.PIPETX07EQCOEFF(pipe_tx07_eq_coeff[17:0])
   ,.PIPETX07EQCONTROL(pipe_tx07_eq_control[1:0])
   ,.PIPETX07EQDEEMPH(pipe_tx07_eq_deemph[5:0])
   ,.PIPETX07EQDONE(pipe_tx07_eq_done)
   ,.PIPETX07POWERDOWN(pipe_tx07_powerdown[1:0])
   ,.PIPETX07STARTBLOCK(pipe_tx07_start_block)
   ,.PIPETX07SYNCHEADER(pipe_tx07_sync_header[1:0])
   ,.PIPETX08CHARISK(pipe_tx08_char_is_k[1:0])
   ,.PIPETX08COMPLIANCE(pipe_tx08_compliance)
   ,.PIPETX08DATA(pipe_tx08_data_out[31:0])
   ,.PIPETX08DATAVALID(pipe_tx08_data_valid)
   ,.PIPETX08ELECIDLE(pipe_tx08_elec_idle)
   ,.PIPETX08EQCOEFF(pipe_tx08_eq_coeff[17:0])
   ,.PIPETX08EQCONTROL(pipe_tx08_eq_control[1:0])
   ,.PIPETX08EQDEEMPH(pipe_tx08_eq_deemph[5:0])
   ,.PIPETX08EQDONE(pipe_tx08_eq_done)
   ,.PIPETX08POWERDOWN(pipe_tx08_powerdown[1:0])
   ,.PIPETX08STARTBLOCK(pipe_tx08_start_block)
   ,.PIPETX08SYNCHEADER(pipe_tx08_sync_header[1:0])
   ,.PIPETX09CHARISK(pipe_tx09_char_is_k[1:0])
   ,.PIPETX09COMPLIANCE(pipe_tx09_compliance)
   ,.PIPETX09DATA(pipe_tx09_data_out[31:0])
   ,.PIPETX09DATAVALID(pipe_tx09_data_valid)
   ,.PIPETX09ELECIDLE(pipe_tx09_elec_idle)
   ,.PIPETX09EQCOEFF(pipe_tx09_eq_coeff[17:0])
   ,.PIPETX09EQCONTROL(pipe_tx09_eq_control[1:0])
   ,.PIPETX09EQDEEMPH(pipe_tx09_eq_deemph[5:0])
   ,.PIPETX09EQDONE(pipe_tx09_eq_done)
   ,.PIPETX09POWERDOWN(pipe_tx09_powerdown[1:0])
   ,.PIPETX09STARTBLOCK(pipe_tx09_start_block)
   ,.PIPETX09SYNCHEADER(pipe_tx09_sync_header[1:0])
   ,.PIPETX10CHARISK(pipe_tx10_char_is_k[1:0])
   ,.PIPETX10COMPLIANCE(pipe_tx10_compliance)
   ,.PIPETX10DATA(pipe_tx10_data_out[31:0])
   ,.PIPETX10DATAVALID(pipe_tx10_data_valid)
   ,.PIPETX10ELECIDLE(pipe_tx10_elec_idle)
   ,.PIPETX10EQCOEFF(pipe_tx10_eq_coeff[17:0])
   ,.PIPETX10EQCONTROL(pipe_tx10_eq_control[1:0])
   ,.PIPETX10EQDEEMPH(pipe_tx10_eq_deemph[5:0])
   ,.PIPETX10EQDONE(pipe_tx10_eq_done)
   ,.PIPETX10POWERDOWN(pipe_tx10_powerdown[1:0])
   ,.PIPETX10STARTBLOCK(pipe_tx10_start_block)
   ,.PIPETX10SYNCHEADER(pipe_tx10_sync_header[1:0])
   ,.PIPETX11CHARISK(pipe_tx11_char_is_k[1:0])
   ,.PIPETX11COMPLIANCE(pipe_tx11_compliance)
   ,.PIPETX11DATA(pipe_tx11_data_out[31:0])
   ,.PIPETX11DATAVALID(pipe_tx11_data_valid)
   ,.PIPETX11ELECIDLE(pipe_tx11_elec_idle)
   ,.PIPETX11EQCOEFF(pipe_tx11_eq_coeff[17:0])
   ,.PIPETX11EQCONTROL(pipe_tx11_eq_control[1:0])
   ,.PIPETX11EQDEEMPH(pipe_tx11_eq_deemph[5:0])
   ,.PIPETX11EQDONE(pipe_tx11_eq_done)
   ,.PIPETX11POWERDOWN(pipe_tx11_powerdown[1:0])
   ,.PIPETX11STARTBLOCK(pipe_tx11_start_block)
   ,.PIPETX11SYNCHEADER(pipe_tx11_sync_header[1:0])
   ,.PIPETX12CHARISK(pipe_tx12_char_is_k[1:0])
   ,.PIPETX12COMPLIANCE(pipe_tx12_compliance)
   ,.PIPETX12DATA(pipe_tx12_data_out[31:0])
   ,.PIPETX12DATAVALID(pipe_tx12_data_valid)
   ,.PIPETX12ELECIDLE(pipe_tx12_elec_idle)
   ,.PIPETX12EQCOEFF(pipe_tx12_eq_coeff[17:0])
   ,.PIPETX12EQCONTROL(pipe_tx12_eq_control[1:0])
   ,.PIPETX12EQDEEMPH(pipe_tx12_eq_deemph[5:0])
   ,.PIPETX12EQDONE(pipe_tx12_eq_done)
   ,.PIPETX12POWERDOWN(pipe_tx12_powerdown[1:0])
   ,.PIPETX12STARTBLOCK(pipe_tx12_start_block)
   ,.PIPETX12SYNCHEADER(pipe_tx12_sync_header[1:0])
   ,.PIPETX13CHARISK(pipe_tx13_char_is_k[1:0])
   ,.PIPETX13COMPLIANCE(pipe_tx13_compliance)
   ,.PIPETX13DATA(pipe_tx13_data_out[31:0])
   ,.PIPETX13DATAVALID(pipe_tx13_data_valid)
   ,.PIPETX13ELECIDLE(pipe_tx13_elec_idle)
   ,.PIPETX13EQCOEFF(pipe_tx13_eq_coeff[17:0])
   ,.PIPETX13EQCONTROL(pipe_tx13_eq_control[1:0])
   ,.PIPETX13EQDEEMPH(pipe_tx13_eq_deemph[5:0])
   ,.PIPETX13EQDONE(pipe_tx13_eq_done)
   ,.PIPETX13POWERDOWN(pipe_tx13_powerdown[1:0])
   ,.PIPETX13STARTBLOCK(pipe_tx13_start_block)
   ,.PIPETX13SYNCHEADER(pipe_tx13_sync_header[1:0])
   ,.PIPETX14CHARISK(pipe_tx14_char_is_k[1:0])
   ,.PIPETX14COMPLIANCE(pipe_tx14_compliance)
   ,.PIPETX14DATA(pipe_tx14_data_out[31:0])
   ,.PIPETX14DATAVALID(pipe_tx14_data_valid)
   ,.PIPETX14ELECIDLE(pipe_tx14_elec_idle)
   ,.PIPETX14EQCOEFF(pipe_tx14_eq_coeff[17:0])
   ,.PIPETX14EQCONTROL(pipe_tx14_eq_control[1:0])
   ,.PIPETX14EQDEEMPH(pipe_tx14_eq_deemph[5:0])
   ,.PIPETX14EQDONE(pipe_tx14_eq_done)
   ,.PIPETX14POWERDOWN(pipe_tx14_powerdown[1:0])
   ,.PIPETX14STARTBLOCK(pipe_tx14_start_block)
   ,.PIPETX14SYNCHEADER(pipe_tx14_sync_header[1:0])
   ,.PIPETX15CHARISK(pipe_tx15_char_is_k[1:0])
   ,.PIPETX15COMPLIANCE(pipe_tx15_compliance)
   ,.PIPETX15DATA(pipe_tx15_data_out[31:0])
   ,.PIPETX15DATAVALID(pipe_tx15_data_valid)
   ,.PIPETX15ELECIDLE(pipe_tx15_elec_idle)
   ,.PIPETX15EQCOEFF(pipe_tx15_eq_coeff[17:0])
   ,.PIPETX15EQCONTROL(pipe_tx15_eq_control[1:0])
   ,.PIPETX15EQDEEMPH(pipe_tx15_eq_deemph[5:0])
   ,.PIPETX15EQDONE(pipe_tx15_eq_done)
   ,.PIPETX15POWERDOWN(pipe_tx15_powerdown[1:0])
   ,.PIPETX15STARTBLOCK(pipe_tx15_start_block)
   ,.PIPETX15SYNCHEADER(pipe_tx15_sync_header[1:0])
   ,.PIPETXDEEMPH(pipe_tx_deemph)
   ,.PIPETXMARGIN(pipe_tx_margin[2:0])
   ,.PIPETXRATE(pipe_tx_rate[1:0])
   ,.PIPETXRCVRDET(pipe_tx_rcvr_det)
   ,.PIPETXRESET(pipe_tx_reset)
   ,.PIPETXSWING(pipe_tx_swing)
   ,.PLEQINPROGRESS(pl_eq_in_progress)
   ,.PLEQPHASE(pl_eq_phase[1:0])
   ,.PLEQRESETEIEOSCOUNT(pl_eq_reset_eieos_count)
   ,.PLGEN2UPSTREAMPREFERDEEMPH(pl_gen2_upstream_prefer_deemph)
   ,.PLGEN34EQMISMATCH(pl_gen34_eq_mismatch)
   ,.PLGEN34REDOEQSPEED(pl_gen34_redo_eq_speed)
   ,.PLGEN34REDOEQUALIZATION(pl_gen34_redo_equalization)
   ,.RESETN(reset_n)
   ,.SAXISCCTDATA(s_axis_cc_tdata_int[255:0])
   ,.SAXISCCTKEEP(s_axis_cc_tkeep_int[7:0])
   ,.SAXISCCTLAST(s_axis_cc_tlast_int)
   ,.SAXISCCTREADY(s_axis_cc_tready_int[3:0])
   ,.SAXISCCTUSER(s_axis_cc_tuser_int[32:0])
   ,.SAXISCCTVALID(s_axis_cc_tvalid_int)
   ,.SAXISRQTDATA(s_axis_rq_tdata_int[255:0])
   ,.SAXISRQTKEEP(s_axis_rq_tkeep_int[7:0])
   ,.SAXISRQTLAST(s_axis_rq_tlast_int)
   ,.SAXISRQTREADY(s_axis_rq_tready_int[3:0])
   ,.SAXISRQTUSER(s_axis_rq_tuser_int[61:0])
   ,.SAXISRQTVALID(s_axis_rq_tvalid_int)
   ,.USERCLK2(user_clk2_to_e4)
   ,.USERCLKEN(user_clk_en_to_e4)
   ,.USERCLK(user_clk_to_e4)
   ,.USERSPAREIN({32{1'b0}})
   ,.USERSPAREOUT( )

  );

  end

  endgenerate

  // BlockRAM Module

  xp4_usp_smsw_bram 
 #(
   .TCQ(TCQ)
  ,.AXISTEN_IF_MSIX_TO_RAM_PIPELINE(AXISTEN_IF_MSIX_TO_RAM_PIPELINE)
  ,.AXISTEN_IF_MSIX_FROM_RAM_PIPELINE(AXISTEN_IF_MSIX_FROM_RAM_PIPELINE)
  ,.TPH_TO_RAM_PIPELINE(TPH_TO_RAM_PIPELINE)
  ,.TPH_FROM_RAM_PIPELINE(TPH_FROM_RAM_PIPELINE)
  ,.TL_COMPLETION_RAM_SIZE(TL_COMPLETION_RAM_SIZE)
  ,.TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE(TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE)
  ,.TL_RX_COMPLETION_TO_RAM_READ_PIPELINE(TL_RX_COMPLETION_TO_RAM_READ_PIPELINE)
  ,.TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE(TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE)
  ,.TL_RX_POSTED_TO_RAM_WRITE_PIPELINE(TL_RX_POSTED_TO_RAM_WRITE_PIPELINE)
  ,.TL_RX_POSTED_TO_RAM_READ_PIPELINE(TL_RX_POSTED_TO_RAM_READ_PIPELINE)
  ,.TL_RX_POSTED_FROM_RAM_READ_PIPELINE(TL_RX_POSTED_FROM_RAM_READ_PIPELINE)
  ,.LL_REPLAY_TO_RAM_PIPELINE(LL_REPLAY_TO_RAM_PIPELINE)
  ,.LL_REPLAY_FROM_RAM_PIPELINE(LL_REPLAY_FROM_RAM_PIPELINE)
  ,.TL_PF_ENABLE_REG(TL_PF_ENABLE_REG)
  ,.SRIOV_CAP_ENABLE(SRIOV_CAP_ENABLE)
  ,.PF0_SRIOV_CAP_TOTAL_VF(PF0_SRIOV_CAP_TOTAL_VF)
  ,.PF1_SRIOV_CAP_TOTAL_VF(PF1_SRIOV_CAP_TOTAL_VF)
  ,.PF2_SRIOV_CAP_TOTAL_VF(PF2_SRIOV_CAP_TOTAL_VF)
  ,.PF3_SRIOV_CAP_TOTAL_VF(PF3_SRIOV_CAP_TOTAL_VF)
  ,.PF0_TPHR_CAP_ENABLE(PF0_TPHR_CAP_ENABLE)
  ,.MSIX_CAP_TABLE_SIZE(MSIX_CAP_TABLE_SIZE)
  ,.MSIX_TABLE_RAM_ENABLE(MSIX_TABLE_RAM_ENABLE)


  ) pcie_4_0_bram_inst (

   .core_clk_i(core_clk)
  ,.user_clk_i(user_clk) 
  ,.reset_i(!reset_n)
  ,.mi_rep_addr_i(mi_replay_ram_address0[8:0])
  ,.mi_rep_wdata_i({mi_replay_ram_write_data1[127:0],mi_replay_ram_write_data0[127:0]})
  ,.mi_rep_wen_i(mi_replay_ram_write_enable0)
  ,.mi_rep_rdata_o({mi_replay_ram_read_data1[127:0],mi_replay_ram_read_data0[127:0]})
  ,.mi_rep_rden_i(mi_replay_ram_read_enable0)
  ,.mi_rep_err_cor_o(mi_replay_ram_err_cor[3:0])
  ,.mi_rep_err_uncor_o(mi_replay_ram_err_uncor[3:0])
  ,.mi_req_waddr0_i(mi_rx_posted_request_ram_write_address0[8:0])
  ,.mi_req_wdata0_i(mi_rx_posted_request_ram_write_data0[143:0])
  ,.mi_req_wen0_i(mi_rx_posted_request_ram_write_enable0)
  ,.mi_req_waddr1_i(mi_rx_posted_request_ram_write_address1[8:0])
  ,.mi_req_wdata1_i(mi_rx_posted_request_ram_write_data1[143:0])
  ,.mi_req_wen1_i(mi_rx_posted_request_ram_write_enable1)
  ,.mi_req_raddr0_i(mi_rx_posted_request_ram_read_address0[8:0])
  ,.mi_req_rdata0_o(mi_rx_posted_request_ram_read_data0[143:0])
  ,.mi_req_ren0_i(mi_rx_posted_request_ram_read_enable0)
  ,.mi_req_raddr1_i(mi_rx_posted_request_ram_read_address1[8:0])
  ,.mi_req_rdata1_o(mi_rx_posted_request_ram_read_data1[143:0])
  ,.mi_req_ren1_i(mi_rx_posted_request_ram_read_enable1)
  ,.mi_req_err_cor_o(mi_rx_posted_request_ram_err_cor[5:0])
  ,.mi_req_err_uncor_o(mi_rx_posted_request_ram_err_uncor[5:0])
  ,.mi_cpl_waddr0_i(mi_rx_completion_ram_write_address0[8:0])
  ,.mi_cpl_wdata0_i(mi_rx_completion_ram_write_data0[143:0])
  ,.mi_cpl_wen0_i(mi_rx_completion_ram_write_enable0[1:0])
  ,.mi_cpl_waddr1_i(mi_rx_completion_ram_write_address1[8:0])
  ,.mi_cpl_wdata1_i(mi_rx_completion_ram_write_data1[143:0])
  ,.mi_cpl_wen1_i(mi_rx_completion_ram_write_enable1[1:0])
  ,.mi_cpl_raddr0_i(mi_rx_completion_ram_read_address0[8:0])
  ,.mi_cpl_rdata0_o(mi_rx_completion_ram_read_data0[143:0])
  ,.mi_cpl_ren0_i(mi_rx_completion_ram_read_enable0[1:0])
  ,.mi_cpl_raddr1_i(mi_rx_completion_ram_read_address1[8:0])
  ,.mi_cpl_rdata1_o(mi_rx_completion_ram_read_data1[143:0])
  ,.mi_cpl_ren1_i(mi_rx_completion_ram_read_enable1[1:0])
  ,.mi_cpl_err_cor_o(mi_rx_completion_ram_err_cor[11:0])
  ,.mi_cpl_err_uncor_o(mi_rx_completion_ram_err_uncor[11:0])
  ,.cfg_msix_waddr_i(cfg_msix_ram_address[12:0])
  ,.cfg_msix_wdata_i(cfg_msix_ram_write_data[31:0])
  ,.cfg_msix_wdip_i(cfg_msix_ram_write_data[35:32])
  ,.cfg_msix_wen_i(cfg_msix_ram_write_byte_enable[3:0])
  ,.cfg_msix_rdata_o(cfg_msix_ram_read_data[31:0])
  ,.cfg_msix_rdop_o(cfg_msix_ram_read_data[35:32])
  ,.cfg_msix_ren_i(cfg_msix_ram_read_enable)
  ,.user_tph_stt_func_num_i(user_tph_stt_func_num[7:0])
  ,.user_tph_stt_index_i(user_tph_stt_index[5:0])
  ,.user_tph_stt_rd_en_i(user_tph_stt_rd_en)
  ,.user_tph_stt_rd_data_o(user_tph_stt_rd_data[7:0])
  ,.cfg_tph_waddr_i(cfg_tph_ram_address[11:0])
  ,.cfg_tph_wdata_i(cfg_tph_ram_write_data[31:0])
  ,.cfg_tph_wdip_i(cfg_tph_ram_write_data[35:32])
  ,.cfg_tph_wen_i(cfg_tph_ram_write_byte_enable[3:0])
  ,.cfg_tph_rdata_o(cfg_tph_ram_read_data[31:0])
  ,.cfg_tph_rdop_o(cfg_tph_ram_read_data[35:32])
  ,.cfg_tph_ren_i(cfg_tph_ram_read_enable)

  );

  assign mi_replay_ram_err_cor[5:4] = 2'b00;
  assign mi_replay_ram_err_uncor[5:4] = 2'b00;

  // Initialization Controller Module

  xp4_usp_smsw_init_ctrl
 #(
    .TCQ(TCQ)
   ,.PL_UPSTREAM_FACING(PL_UPSTREAM_FACING)
   ,.IS_SWITCH_PORT(IS_SWITCH_PORT)
   ,.CRM_CORE_CLK_FREQ_500(CRM_CORE_CLK_FREQ_500)
   ,.CRM_USER_CLK_FREQ(CRM_USER_CLK_FREQ)

  ) pcie_4_0_init_ctrl_inst ( 

    .core_clk_i (core_clk)
   ,.user_clk_i (user_clk)
   ,.reset_n_o (reset_n)
   ,.pipe_reset_n_o (pipe_reset_n)
   ,.mgmt_reset_n_o (mgmt_reset_n)
   ,.mgmt_sticky_reset_n_o (mgmt_sticky_reset_n)
   ,.phy_rdy_i (phy_rdy)
   ,.cfg_hot_reset_in_i(cfg_hot_reset_in)
   ,.cfg_phy_link_down_i(cfg_phy_link_down_wire)
   ,.cfg_phy_link_down_user_clk_o(cfg_phy_link_down_user_clk)
   ,.state_o ()
   ,.user_clk_en_o(user_clk_en)
   ,.user_clkgate_en_o(user_clkgate_en)

  );

  // VF Decode Module
  
  xp4_usp_smsw_vf_decode
 #(
    .TCQ(TCQ)
   ,.TL_PF_ENABLE_REG(TL_PF_ENABLE_REG)
   ,.PF0_SRIOV_CAP_TOTAL_VF(PF0_SRIOV_CAP_TOTAL_VF)
   ,.PF1_SRIOV_CAP_TOTAL_VF(PF1_SRIOV_CAP_TOTAL_VF)
   ,.PF2_SRIOV_CAP_TOTAL_VF(PF2_SRIOV_CAP_TOTAL_VF)
   ,.PF3_SRIOV_CAP_TOTAL_VF(PF3_SRIOV_CAP_TOTAL_VF)
   ,.PF0_SRIOV_FIRST_VF_OFFSET(PF0_SRIOV_FIRST_VF_OFFSET)
   ,.PF1_SRIOV_FIRST_VF_OFFSET(PF1_SRIOV_FIRST_VF_OFFSET)
   ,.PF2_SRIOV_FIRST_VF_OFFSET(PF2_SRIOV_FIRST_VF_OFFSET)
   ,.PF3_SRIOV_FIRST_VF_OFFSET(PF3_SRIOV_FIRST_VF_OFFSET)
   ,.SRIOV_CAP_ENABLE(SRIOV_CAP_ENABLE)
   ,.ARI_CAP_ENABLE(ARI_CAP_ENABLE)

  ) pcie_4_0_vf_decode_inst (

     .clk_i(user_clk)
    ,.reset_i(!reset_n)
    ,.link_down_i(cfg_phy_link_down_user_clk)
    ,.cfg_ext_write_received_i(cfg_ext_write_received)
    ,.cfg_ext_register_number_i(cfg_ext_register_number[9:0])
    ,.cfg_ext_function_number_i(cfg_ext_function_number[7:0])
    ,.cfg_ext_write_data_i(cfg_ext_write_data[31:0])
    ,.cfg_ext_write_byte_enable_i(cfg_ext_write_byte_enable[3:0])
    ,.cfg_flr_in_process_i(cfg_flr_in_process[3:0])

    ,.cfg_vf_flr_in_process_o(cfg_vf_flr_in_process[251:0])
    ,.cfg_vf_status_o(cfg_vf_status[503:0])
    ,.cfg_vf_power_state_o(cfg_vf_power_state[755:0])
    ,.cfg_vf_tph_requester_enable_o(cfg_vf_tph_requester_enable[251:0])
    ,.cfg_vf_tph_st_mode_o(cfg_vf_tph_st_mode[755:0])
    ,.cfg_interrupt_msix_vf_enable_o(cfg_interrupt_msix_vf_enable[251:0])
    ,.cfg_interrupt_msix_vf_mask_o(cfg_interrupt_msix_vf_mask[251:0])

  );

  // PL EQ Interface Module

  xp4_usp_smsw_pl_eq
 #(
     .TCQ(TCQ)
    ,.IMPL_TARGET(IMPL_TARGET)
    ,.PL_UPSTREAM_FACING(PL_UPSTREAM_FACING)

  ) pcie_4_0_pl_eq_inst (

     .clk_i(user_clk)
    ,.reset_i(!reset_n)
    ,.link_down_reset_i(cfg_phy_link_down_user_clk)

    ,.cfg_ltssm_state_i(cfg_ltssm_state[5:0])     
    ,.pl_redo_eq_i(pl_redo_eq)
    ,.pl_redo_eq_speed_i(pl_redo_eq_speed)
    ,.pl_eq_mismatch_o(pl_eq_mismatch)
    ,.pl_redo_eq_pending_o(pl_redo_eq_pending)
    ,.pl_gen34_redo_equalization_o(pl_gen34_redo_equalization)
    ,.pl_gen34_redo_eq_speed_o(pl_gen34_redo_eq_speed)
    ,.pl_gen34_eq_mismatch_i(pl_gen34_eq_mismatch)

  );

  // AXI4ST 256b/512b Bridge Module
  xp4_usp_smsw_512b_intfc
 #(
        .TCQ(TCQ),
        .IMPL_TARGET(IMPL_TARGET),
        .AXISTEN_IF_EXT_512_INTFC_RAM_STYLE(AXISTEN_IF_EXT_512_INTFC_RAM_STYLE),
        .AXI4_USER_DATA_WIDTH(AXI4_DATA_WIDTH),
        .AXI4_CORE_DATA_WIDTH(256),
        .AXI4_USER_CQ_TUSER_WIDTH(AXI4_CQ_TUSER_WIDTH),
        .AXI4_USER_CC_TUSER_WIDTH(AXI4_CC_TUSER_WIDTH),
        .AXI4_USER_RQ_TUSER_WIDTH(AXI4_RQ_TUSER_WIDTH),
        .AXI4_USER_RC_TUSER_WIDTH(AXI4_RC_TUSER_WIDTH),
        .AXI4_CORE_CQ_TUSER_WIDTH(88),
        .AXI4_CORE_CC_TUSER_WIDTH(33),
        .AXI4_CORE_RQ_TUSER_WIDTH(62),
        .AXI4_CORE_RC_TUSER_WIDTH(75),
        .AXI4_USER_CQ_TKEEP_WIDTH(AXI4_TKEEP_WIDTH),
        .AXI4_USER_CC_TKEEP_WIDTH(AXI4_TKEEP_WIDTH),
        .AXI4_USER_RQ_TKEEP_WIDTH(AXI4_TKEEP_WIDTH),
        .AXI4_USER_RC_TKEEP_WIDTH(AXI4_TKEEP_WIDTH),
        .AXI4_CORE_CQ_TKEEP_WIDTH(8),
        .AXI4_CORE_CC_TKEEP_WIDTH(8),
        .AXI4_CORE_RQ_TKEEP_WIDTH(8),
        .AXI4_CORE_RC_TKEEP_WIDTH(8),
        .AXI4_CORE_CQ_TREADY_WIDTH(22),
        .AXI4_CORE_RC_TREADY_WIDTH(22),

        .AXISTEN_IF_EXT_512_CQ_STRADDLE(AXISTEN_IF_EXT_512_CQ_STRADDLE),
        .AXISTEN_IF_EXT_512_CC_STRADDLE(AXISTEN_IF_EXT_512_CC_STRADDLE),
        .AXISTEN_IF_EXT_512_RQ_STRADDLE(AXISTEN_IF_EXT_512_RQ_STRADDLE),
        .AXISTEN_IF_EXT_512_RC_STRADDLE(AXISTEN_IF_EXT_512_RC_STRADDLE),
        .AXISTEN_IF_EXT_512_RC_4TLP_STRADDLE(AXISTEN_IF_EXT_512_RC_4TLP_STRADDLE),
        .AXISTEN_IF_CQ_ALIGNMENT_MODE(AXISTEN_IF_CQ_ALIGNMENT_MODE),
        .AXISTEN_IF_CC_ALIGNMENT_MODE(AXISTEN_IF_CC_ALIGNMENT_MODE),
        .AXISTEN_IF_RQ_ALIGNMENT_MODE(AXISTEN_IF_RQ_ALIGNMENT_MODE),
        .AXISTEN_IF_RC_ALIGNMENT_MODE(AXISTEN_IF_RC_ALIGNMENT_MODE),
        .AXISTEN_IF_RQ_CC_REGISTERED_TREADY(AXISTEN_IF_RQ_CC_REGISTERED_TREADY),
        .AXISTEN_IF_RX_PARITY_EN(AXISTEN_IF_RX_PARITY_EN),
        .AXISTEN_IF_TX_PARITY_EN(AXISTEN_IF_TX_PARITY_EN)

     ) pcie4_0_512b_intfc_mod (

        .user_clk_i         (user_clk),
        .user_clk2_i        (user_clk2),
        .user_clk_en_i      (user_clk_en),
        .reset_n_user_clk_i (reset_n),
        .reset_n_user_clk2_i(reset_n),
        .link_down_reset_i  (cfg_phy_link_down_user_clk),
        //-----------------------------------
        // Client-side signals
        //-----------------------------------
        // CQ Interface
        .m_axis_cq_tdata_o  (m_axis_cq_tdata),
        .m_axis_cq_tvalid_o (m_axis_cq_tvalid),
        .m_axis_cq_tuser_o  (m_axis_cq_tuser),
        .m_axis_cq_tlast_o  (m_axis_cq_tlast),
        .m_axis_cq_tkeep_o  (m_axis_cq_tkeep),
        .m_axis_cq_tready_i (m_axis_cq_tready[0]),
        .pcie_cq_np_req_i   (pcie_cq_np_req),
        .pcie_cq_np_req_count_o(pcie_cq_np_req_count_axi512),
        // CC Interface
        .s_axis_cc_tdata_i  (s_axis_cc_tdata),
        .s_axis_cc_tvalid_i (s_axis_cc_tvalid),
        .s_axis_cc_tuser_i  (s_axis_cc_tuser),
        .s_axis_cc_tlast_i  (s_axis_cc_tlast),
        .s_axis_cc_tkeep_i  (s_axis_cc_tkeep),
        .s_axis_cc_tready_o (s_axis_cc_tready_axi512),
        // RQ Interface
        .s_axis_rq_tdata_i  (s_axis_rq_tdata),
        .s_axis_rq_tvalid_i (s_axis_rq_tvalid),
        .s_axis_rq_tuser_i  (s_axis_rq_tuser),
        .s_axis_rq_tlast_i  (s_axis_rq_tlast),
        .s_axis_rq_tkeep_i  (s_axis_rq_tkeep),
        .s_axis_rq_tready_o (s_axis_rq_tready_axi512),
        // RC Interface
        .m_axis_rc_tdata_o  (m_axis_rc_tdata),
        .m_axis_rc_tvalid_o (m_axis_rc_tvalid),
        .m_axis_rc_tuser_o  (m_axis_rc_tuser),
        .m_axis_rc_tlast_o  (m_axis_rc_tlast),
        .m_axis_rc_tkeep_o  (m_axis_rc_tkeep),
        .m_axis_rc_tready_i (m_axis_rc_tready[0]),
        //-----------------------------------
        // Core-side signals
        //-----------------------------------
        // CQ Interface
        .core_cq_tdata_i    (m_axis_cq_tdata_int),
        .core_cq_tvalid_i   (m_axis_cq_tvalid_int),
        .core_cq_tuser_i    (m_axis_cq_tuser_int),
        .core_cq_tlast_i    (m_axis_cq_tlast_int),
        .core_cq_tkeep_i    (m_axis_cq_tkeep_int),
        .core_cq_tready_o   (m_axis_cq_tready_axi512),
        .posted_req_delivered_o(pcie_posted_req_delivered),
        .cq_pipeline_empty_o(pcie_cq_pipeline_empty),
        .cq_np_user_credit_rcvd_o(pcie_cq_np_user_credit_rcvd),
        // CC Interface
        .core_cc_tdata_o    (s_axis_cc_tdata_axi512),
        .core_cc_tvalid_o   (s_axis_cc_tvalid_axi512),
        .core_cc_tuser_o    (s_axis_cc_tuser_axi512),
        .core_cc_tlast_o    (s_axis_cc_tlast_axi512),
        .core_cc_tkeep_o    (s_axis_cc_tkeep_axi512),
        .core_cc_tready_i   (s_axis_cc_tready_int),
        // RQ Interface
        .core_rq_tdata_o    (s_axis_rq_tdata_axi512),
        .core_rq_tvalid_o   (s_axis_rq_tvalid_axi512),
        .core_rq_tuser_o    (s_axis_rq_tuser_axi512),
        .core_rq_tlast_o    (s_axis_rq_tlast_axi512),
        .core_rq_tkeep_o    (s_axis_rq_tkeep_axi512),
        .core_rq_tready_i   (s_axis_rq_tready_int),
        // RC Interface
        .core_rc_tdata_i    (m_axis_rc_tdata_int),
        .core_rc_tvalid_i   (m_axis_rc_tvalid_int),
        .core_rc_tuser_i    (m_axis_rc_tuser_int),
        .core_rc_tlast_i    (m_axis_rc_tlast_int),
        .core_rc_tkeep_i    (m_axis_rc_tkeep_int),
        .core_rc_tready_o   (m_axis_rc_tready_axi512),
        .compl_delivered_o  (pcie_compl_delivered),
        .compl_delivered_tag0_o(pcie_compl_delivered_tag0),
        .compl_delivered_tag1_o(pcie_compl_delivered_tag1)
        );

      assign s_axis_cc_tdata_int = s_axis_cc_tdata_axi512;
      assign s_axis_cc_tvalid_int = s_axis_cc_tvalid_axi512;
      assign s_axis_cc_tuser_int = s_axis_cc_tuser_axi512;
      assign s_axis_cc_tlast_int = s_axis_cc_tlast_axi512;
      assign s_axis_cc_tkeep_int = s_axis_cc_tkeep_axi512;
      
      assign s_axis_rq_tdata_int = s_axis_rq_tdata_axi512;
      assign s_axis_rq_tvalid_int = s_axis_rq_tvalid_axi512;
      assign s_axis_rq_tuser_int = s_axis_rq_tuser_axi512;
      assign s_axis_rq_tlast_int = s_axis_rq_tlast_axi512;
      assign s_axis_rq_tkeep_int = s_axis_rq_tkeep_axi512;

    
   assign m_axis_cq_tready_int[21:0] = (AXISTEN_IF_EXT_512 == "TRUE") ? 
                                                           m_axis_cq_tready_axi512 :
                                                           m_axis_cq_tready;

   assign m_axis_rc_tready_int[21:0] = (AXISTEN_IF_EXT_512 == "TRUE") ? 
                                                           m_axis_rc_tready_axi512 :
                                                           m_axis_rc_tready;

   assign s_axis_cc_tready = (AXISTEN_IF_EXT_512 == "TRUE") ? {4{s_axis_cc_tready_axi512}} :
                                                              s_axis_cc_tready_int;

   assign s_axis_rq_tready = (AXISTEN_IF_EXT_512 == "TRUE") ? {4{s_axis_rq_tready_axi512}} :
                                                              s_axis_rq_tready_int;

   assign pcie_cq_np_req_count = (AXISTEN_IF_EXT_512 == "TRUE") ? pcie_cq_np_req_count_axi512:
                                                                  pcie_cq_np_req_count_int;

  generate if ((TL_USER_SPARE[1]) ||
               ((CRM_CORE_CLK_FREQ_500 == "TRUE") && (CRM_USER_CLK_FREQ[1:0] == 2'b11)) ||
               ((CRM_CORE_CLK_FREQ_500 == "FALSE") && (CRM_USER_CLK_FREQ[1:0] == 2'b10))) begin: seqnum_fifo_bypass
  
    assign pcie_rq_seq_num0[5:0] = pcie_rq_seq_num0_cc[5:0];
    assign pcie_rq_seq_num_vld0 = pcie_rq_seq_num_vld0_cc;
  
  end else begin: seqnum_fifo
  
     //
     // Sequence Number FIFOs
     //

  xp4_usp_smsw_seqnum_fifo #(
     .RAM_WIDTH(7), 
     .RAM_DEPTH(16), 
     .FIFO_FULL_HIGH_THRESHOLD(16),
     .ADDR_WIDTH(4)
   ) seq_fifo_0 (
     .core_reset_n_i(reset_n),
     .core_clk_i(core_clk),
     .user_reset_n_i(reset_n),
     .user_clk_i(user_clk),
     .data_i({pcie_rq_seq_num_vld0_cc, pcie_rq_seq_num0_cc[5:0]}),
     .data_o({pcie_rq_seq_num_vld0, pcie_rq_seq_num0[5:0]})
   );

  end
  endgenerate


endmodule

//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_init_ctrl.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
//**  Description: PCI Express Gen4 Block Initialization Controller
//**  Revision: $Revision: #19 $
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_init_ctrl #(
     parameter           TCQ = 100
   , parameter           PL_UPSTREAM_FACING = "TRUE"
   , parameter           IS_SWITCH_PORT = "FALSE"
   , parameter           CRM_CORE_CLK_FREQ_500="TRUE"
   , parameter [1:0]     CRM_USER_CLK_FREQ=2'b10
)(
  input  wire         core_clk_i,
  input  wire         user_clk_i,
  input  wire         phy_rdy_i,
  input  wire         cfg_hot_reset_in_i,
  input  wire         cfg_phy_link_down_i,
  output reg          cfg_phy_link_down_user_clk_o,
  output wire   [2:0] state_o,

  (* keep = "true", max_fanout = 1000 *) output reg          reset_n_o,
  output wire                                                pipe_reset_n_o,
  (* keep = "true", max_fanout = 1000 *) output reg          mgmt_reset_n_o,
  (* keep = "true", max_fanout = 1000 *) output reg          mgmt_sticky_reset_n_o,

  output wire         user_clk_en_o,
  output wire         user_clkgate_en_o
  );

   localparam STATE_RESET   = 3'b000;
   localparam STATE_MGMT_RESET_DEASSERT = 3'b001;
   localparam STATE_PHY_RDY = 3'b100;
   localparam STATE_RESET_DEASSERT = 3'b101;
   
   localparam CLK_QUARTER0  = 3'b0_00; // core=250, user=62.5, user2 = 62.5 
   localparam CLK_HALF0     = 3'b0_01; // core=250, user=125,  user2 = 125
   localparam CLK_EQUAL0    = 3'b0_10; // core=250, user=250,  user2 = 250
   localparam CLK_INVALID0  = 3'b0_11; // core=250, user=250,  user2 = 500
   localparam CLK_INVALID1  = 3'b1_00; // core=500, user=62.5, user2 = 62.5
   localparam CLK_QUARTER1  = 3'b1_01; // core=500, user=125,  user2 = 125
   localparam CLK_HALF1     = 3'b1_10; // core=500, user=250,  user2 = 250
   localparam CLK_HALF2     = 3'b1_11; // core=500, user=250,  user2 = 500

   reg           [2:0] reg_state;
   reg           [2:0] reg_next_state;
   reg           [1:0] reg_phy_rdy = 2'b11;
   reg           [1:0] reg_cold_reset = 2'b11;
   reg                 reg_reset_n_o;
   reg                 reg_pipe_reset_n_o;
   reg                 reg_mgmt_reset_n_o;
   reg                 reg_mgmt_sticky_reset_n_o;
   reg           [1:0] reg_reset_timer;
   wire          [2:0] state_w;
   wire          [2:0] next_state_w;
   wire                phy_rdy;
   wire                cold_reset_n;
   wire          [1:0] reset_timer_w;
   wire                attr_pl_upstream_facing;
   wire                attr_is_switch_port;

   wire 	       attr_crm_core_clk_freq_500;
   wire [1:0] 	       attr_crm_user_clk_freq;
   wire 	       user2_eq_core;
   reg [1:0] 	       counter;
   
   (* keep = "true", max_fanout = 1000 *) reg 		       user_clk_en_int;
   
   reg 		       user_clkgate_en_int;
   
   
   assign attr_crm_core_clk_freq_500 = (CRM_CORE_CLK_FREQ_500 == "TRUE") ? 1'b1 : 1'b0;
   assign attr_crm_user_clk_freq = CRM_USER_CLK_FREQ[1:0];
				       
   wire [2:0]  coreuser_clk_ratio  = {attr_crm_core_clk_freq_500, attr_crm_user_clk_freq};

  // common values for {attr_crm_core_clk_freq_500, attr_crm_user_clk_freq}
  // attr_crm_core_clk_freq_500,
  // 0 == 250, 1 == 500
  // attr_crm_user_clk_freq,
  // 0 = 62.5/62.5, 1 = 125/125, 2 = 250/250, 3 = 250/500
  //---------------------------------------------------
  // ratios: c:u(:u2)
  // 0/0 250:62.5(62.5)  -> 1/4(/4) CLK_QUARTER0       // user2_eq_core == 0
  // 0/1 250:125 (125)   -> 1/2(/2) CLK_HALF0          // user2_eq_core == 0
  // 0/2 250:250 (250)   -> 1/1(/1) CLK_EQUAL0         // user2_eq_core == 0
  // 0/3 250:250 (500)   -> 1/1(x2) CLK_INVALID0/EQUAL // user2_eq_core == 1
  // 1/0 500:62.5(62.5)  -> 1/8(/8) CLK_INVALID1/EQUAL // user2_eq_core == 0
  // 1/1 500:125 (125)   -> 1/4(/4) CLK_QUARTER1       // user2_eq_core == 0
  // 1/2 500:250 (250)   -> 1/2(/2) CLK_HALF1          // user2_eq_core == 0
  // 1/3 500:250 (500)   -> 1/2(/1) CLK_HALF2          // user2_eq_core == 1
   
   // user2_eq_core high when user_clk2 is equal to core_clk (and faster than user_clk) else equal to user_clk
   //OBSOLETE// assign user2_eq_core = {attr_crm_user_clk_freq == 2'b11};
      
   // when user2_clk is same as core_clk assign coreuser2_clk_ratio to EQUAL, else
   // user2_clk is same as user_clk so use the coreuser_clk_ratio
   //OBSOLETE// wire [2:0]  coreuser2_clk_ratio = user2_eq_core ? CLK_EQUAL0 : coreuser_clk_ratio;


  always @(posedge core_clk_i or negedge mgmt_reset_n_o) begin

    // hold the count during power-on reset
    if (!mgmt_reset_n_o) begin
      user_clkgate_en_int  <= #TCQ 1'b0;
      user_clk_en_int      <= #TCQ 1'b0;
      counter              <= #TCQ 2'h0;
    // normal free-running operation
    end else begin
      // counter always increments and rolls over, no matter the ratio
      counter <= #TCQ counter + 1;

      // Choose the valid based on the table above
      case (coreuser_clk_ratio)
        CLK_HALF0, CLK_HALF1, CLK_HALF2: begin
	   // one core_clk cycle advanced for _e4 input
          user_clkgate_en_int <= #TCQ counter[0];
          user_clk_en_int     <= #TCQ !counter[0];
        end
        CLK_QUARTER0, CLK_QUARTER1: begin
	   // one core_clk cycle advanced for _e4 input 
          user_clkgate_en_int <= #TCQ (counter == 2'h1);
          user_clk_en_int     <= #TCQ (counter == 2'h2);
        end
        default: begin  // and CLK_EQUAL* case which ties off to high
          user_clkgate_en_int <= #TCQ 1'b1;
          user_clk_en_int     <= #TCQ 1'b1;
        end
      endcase

    end

  end
  // user_clk_en generation
 
  assign attr_pl_upstream_facing = (PL_UPSTREAM_FACING == "TRUE") ? 1'b1 : 1'b0 ;
  assign attr_is_switch_port     = (IS_SWITCH_PORT == "TRUE") ? 1'b1 : 1'b0 ;

  // Generate PHY Ready

  always @(posedge user_clk_i or negedge phy_rdy_i)
  begin
    if (!phy_rdy_i)
      reg_phy_rdy[1:0] <= #TCQ 2'b11;
    else
      reg_phy_rdy[1:0] <= #TCQ {reg_phy_rdy[0], 1'b0};
  end

  assign phy_rdy = !reg_phy_rdy[1];
  
   // Generate Cold reset

  always @(posedge user_clk_i)
  begin
    if (!phy_rdy && reg_cold_reset[1] )
      reg_cold_reset[1:0] <= #TCQ 2'b11;
    else
      reg_cold_reset[1:0] <= #TCQ {reg_cold_reset[0], 1'b0};
  end

  assign cold_reset_n = !reg_cold_reset[1];
  
  // Reset Timer
  
  always @(posedge user_clk_i or negedge phy_rdy_i)
  begin
    if (!phy_rdy_i)
        reg_reset_timer <= #TCQ 2'b00;
    else if ((state_w == STATE_MGMT_RESET_DEASSERT) && (reset_timer_w != 2'b11))
        reg_reset_timer <= #TCQ reset_timer_w + 1'b1;
    else
        reg_reset_timer <= #TCQ reset_timer_w;    
  end
  
  
  // Reset SM
  
  always @(posedge user_clk_i or negedge cold_reset_n)
  begin
    if (!cold_reset_n)
      reg_state <= #TCQ STATE_RESET;
    else
      reg_state <= #TCQ reg_next_state;
  end
  
  always @* begin

    if (attr_pl_upstream_facing) begin // Design is a Upstream Port 

      reg_next_state = STATE_RESET;
      reg_mgmt_reset_n_o = 1'b1;
      reg_mgmt_sticky_reset_n_o = 1'b1;
      reg_reset_n_o = 1'b0;
      reg_pipe_reset_n_o = 1'b0;
      case (state_w)
        STATE_RESET:
        begin
          reg_mgmt_reset_n_o = 1'b0;
          reg_mgmt_sticky_reset_n_o = 1'b0;
          if (phy_rdy)
            reg_next_state = STATE_MGMT_RESET_DEASSERT;
          else
            reg_next_state = STATE_RESET;
          end
        STATE_MGMT_RESET_DEASSERT:
        begin
          if (reset_timer_w == 2'b11)
          reg_next_state = STATE_RESET_DEASSERT;
          else
          reg_next_state = STATE_MGMT_RESET_DEASSERT;
        end
        STATE_RESET_DEASSERT:
        begin
          reg_reset_n_o = 1'b1;
          reg_pipe_reset_n_o = 1'b1;
          if (!phy_rdy)
            reg_next_state = STATE_RESET;
          else
            reg_next_state = STATE_RESET_DEASSERT;
            end
      endcase

    end else  begin // Design is a Downstream Port
      
      reg_next_state = STATE_RESET;
      reg_mgmt_reset_n_o = 1'b1;
      reg_mgmt_sticky_reset_n_o = 1'b1;
      reg_reset_n_o = 1'b0;
      reg_pipe_reset_n_o = 1'b0;
      case (state_w)
        STATE_RESET:
        begin
          reg_mgmt_reset_n_o = 1'b0;
          reg_mgmt_sticky_reset_n_o = 1'b0;
          if (phy_rdy)
            reg_next_state = STATE_MGMT_RESET_DEASSERT;
          else
            reg_next_state = STATE_RESET;
        end
        STATE_MGMT_RESET_DEASSERT:
        begin
          if (reset_timer_w == 2'b11)
            reg_next_state = STATE_PHY_RDY;
          else
            reg_next_state = STATE_MGMT_RESET_DEASSERT;
          end
        STATE_PHY_RDY:
        begin
          if (phy_rdy)
            reg_next_state = STATE_RESET_DEASSERT;
          else
            reg_next_state = STATE_PHY_RDY;
        end
        STATE_RESET_DEASSERT:
        begin
          reg_reset_n_o = 1'b1;
          reg_pipe_reset_n_o = 1'b1;
          if (!phy_rdy)
            reg_next_state = STATE_PHY_RDY;
          else if (attr_is_switch_port && cfg_hot_reset_in_i) begin  // Downstream Port Only
            reg_next_state = STATE_RESET_DEASSERT;
            reg_mgmt_reset_n_o = 1'b0;  
          end else
            reg_next_state = STATE_RESET_DEASSERT;
        end
      endcase
     
    end

  end // 

  // Reset registers pipeline

  (* keep = "true", max_fanout = 1000 *) reg reg_reset_n_2;
  (* keep = "true", max_fanout = 1000 *) reg mgmt_reset_n_2;
  (* keep = "true", max_fanout = 1000 *) reg mgmt_sticky_reset_n_2;
  
  always @(posedge user_clk_i or negedge phy_rdy)
  begin
    if (!phy_rdy)
    begin
      reg_reset_n_2         <= #TCQ 1'b0;
      mgmt_reset_n_2        <= #TCQ 1'b0;
      mgmt_sticky_reset_n_2 <= #TCQ 1'b0;
      
      reset_n_o             <= #TCQ 1'b0;
      mgmt_reset_n_o        <= #TCQ 1'b0;
      mgmt_sticky_reset_n_o <= #TCQ 1'b0;
    end
    else
    begin
      reg_reset_n_2         <= #TCQ reg_reset_n_o;
      mgmt_reset_n_2        <= #TCQ reg_mgmt_reset_n_o;
      mgmt_sticky_reset_n_2 <= #TCQ reg_mgmt_sticky_reset_n_o;
      
      reset_n_o             <= #TCQ reg_reset_n_2;
      mgmt_reset_n_o        <= #TCQ mgmt_reset_n_2;
      mgmt_sticky_reset_n_o <= #TCQ mgmt_sticky_reset_n_2;
    end
  end

   assign state_w = reg_state;
   assign next_state_w = reg_next_state;
   assign pipe_reset_n_o = reg_pipe_reset_n_o;
   assign state_o = reg_state;
   assign reset_timer_w = reg_reset_timer;

   assign user_clkgate_en_o  = user_clkgate_en_int;

   assign user_clk_en_o  = user_clk_en_int;

     // Retime cfg_phy_link_down to user clock

  always @(posedge user_clk_i or negedge phy_rdy)
  begin
    if (!phy_rdy)
      cfg_phy_link_down_user_clk_o <= #TCQ 1'b1;
    else
      cfg_phy_link_down_user_clk_o <= #TCQ cfg_phy_link_down_i;
  end

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_phy_ff_chain.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
/*****************************************************************************
** Description:
**    Flop Chain
**
******************************************************************************/

`timescale 1ps/1ps

`define AS_PHYREG(clk, reset, q, d, rstval)  \
   always @(posedge clk or posedge reset) begin \
      if (reset) \
         q  <= #(TCQ)   rstval;  \
      else  \
         q  <= #(TCQ)   d; \
   end

`define PHYREG(clk, reset, q, d, rstval)  \
   always @(posedge clk) begin \
      if (reset) \
         q  <= #(TCQ)   rstval;  \
      else  \
         q  <= #(TCQ)   d; \
   end

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_phy_ff_chain #(
   // Parameters
   parameter integer PIPELINE_STAGES   = 0,        // 0 = no pipeline; 1 = 1 stage; 2 = 2 stages; 3 = 3 stages
   parameter         ASYNC             = "FALSE",
   parameter integer FF_WIDTH          = 1,
   parameter integer RST_VAL           = 0,
   parameter integer TCQ               = 1
)  (   
   input  wire                         clock_i,          
   input  wire                         reset_i,           
   input  wire [FF_WIDTH-1:0]          ff_i,            
   output wire [FF_WIDTH-1:0]          ff_o        
   );

   genvar   var_i;

   reg   [FF_WIDTH-1:0]          ff_chain [PIPELINE_STAGES:0];

   always @(*) ff_chain[0] = ff_i;

generate
   if (PIPELINE_STAGES > 0) begin:  with_ff_chain
      for (var_i = 0; var_i < PIPELINE_STAGES; var_i = var_i + 1) begin: ff_chain_gen
         if (ASYNC == "TRUE") begin: async_rst
            `AS_PHYREG(clock_i, reset_i, ff_chain[var_i+1], ff_chain[var_i], RST_VAL)
         end else begin: sync_rst
            `PHYREG(clock_i, reset_i, ff_chain[var_i+1], ff_chain[var_i], RST_VAL)
         end
      end
   end
endgenerate

   assign ff_o = ff_chain[PIPELINE_STAGES];

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_phy_pipeline.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
/*****************************************************************************
** Description:
**    Programmable stages for routing to PHY Lanes
**
******************************************************************************/

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_phy_pipeline #(
   // Parameters
   parameter integer PIPELINE_STAGES   = 0,        // 0 = no pipeline; 1 = 1 stage; 2 = 2 stages; 3 = 3 stages
   parameter integer PHY_LANE          = 1,        // Valid settings: 1, 2, 4, 8, 16(only for Gen1/2/3)
   parameter integer TCQ               = 1
)  (   
   // Clock & Reset
   input  wire                         phy_pclk,          
   input  wire                         phy_rst,           
  
   // TX Data 
   input  wire [(PHY_LANE*64)-1:0]     phy_txdata_i,            
   input  wire [(PHY_LANE* 2)-1:0]     phy_txdatak_i,    
   input  wire [PHY_LANE-1:0]          phy_txdata_valid_i,
   input  wire [PHY_LANE-1:0]          phy_txstart_block_i,      
   input  wire [(PHY_LANE* 2)-1:0]     phy_txsync_header_i,      

   output wire [(PHY_LANE*64)-1:0]     phy_txdata_o,            
   output wire [(PHY_LANE* 2)-1:0]     phy_txdatak_o,    
   output wire [PHY_LANE-1:0]          phy_txdata_valid_o,
   output wire [PHY_LANE-1:0]          phy_txstart_block_o,      
   output wire [(PHY_LANE* 2)-1:0]     phy_txsync_header_o,     

   // RX Data
   input  wire [(PHY_LANE*64)-1:0]     phy_rxdata_i,            
   input  wire [(PHY_LANE* 2)-1:0]     phy_rxdatak_i,       
   input  wire [PHY_LANE-1:0]          phy_rxdata_valid_i,         
   input  wire [(PHY_LANE* 2)-1:0]     phy_rxstart_block_i,        
   input  wire [(PHY_LANE* 2)-1:0]     phy_rxsync_header_i,        

   output wire [(PHY_LANE*64)-1:0]     phy_rxdata_o,            
   output wire [(PHY_LANE* 2)-1:0]     phy_rxdatak_o,       
   output wire [PHY_LANE-1:0]          phy_rxdata_valid_o,         
   output wire [(PHY_LANE* 2)-1:0]     phy_rxstart_block_o,        
   output wire [(PHY_LANE* 2)-1:0]     phy_rxsync_header_o,        

   // PHY Command
   input  wire                         phy_txdetectrx_i,        
   input  wire [PHY_LANE-1:0]          phy_txelecidle_i,        
   input  wire [PHY_LANE-1:0]          phy_txcompliance_i,      
   input  wire [PHY_LANE-1:0]          phy_rxpolarity_i,        
   input  wire [1:0]                   phy_powerdown_i,         
   input  wire [1:0]                   phy_rate_i,  

   output wire                         phy_txdetectrx_o,        
   output wire [PHY_LANE-1:0]          phy_txelecidle_o,        
   output wire [PHY_LANE-1:0]          phy_txcompliance_o,      
   output wire [PHY_LANE-1:0]          phy_rxpolarity_o,        
   output wire [1:0]                   phy_powerdown_o,         
   output wire [1:0]                   phy_rate_o,              
    
   // PHY Status
   input  wire [PHY_LANE-1:0]          phy_rxvalid_i,               
   input  wire [PHY_LANE-1:0]          phy_phystatus_i,          
   input  wire [PHY_LANE-1:0]          phy_rxelecidle_i,         
   input  wire [(PHY_LANE*3)-1:0]      phy_rxstatus_i,   

   output wire [PHY_LANE-1:0]          phy_rxvalid_o,               
   output wire [PHY_LANE-1:0]          phy_phystatus_o,          
   output wire [PHY_LANE-1:0]          phy_rxelecidle_o,         
   output wire [(PHY_LANE*3)-1:0]      phy_rxstatus_o,   

   // TX Driver
   input  wire [ 2:0]                  phy_txmargin_i,          
   input  wire                         phy_txswing_i,           
   input  wire                         phy_txdeemph_i,  

   output wire [ 2:0]                  phy_txmargin_o,          
   output wire                         phy_txswing_o,           
   output wire                         phy_txdeemph_o,    
    
   // TX Equalization (Gen3/4)
   input  wire [(PHY_LANE*2)-1:0]      phy_txeq_ctrl_i,      
   input  wire [(PHY_LANE*4)-1:0]      phy_txeq_preset_i,       
   input  wire [(PHY_LANE*6)-1:0]      phy_txeq_coeff_i,   

   output wire [(PHY_LANE*2)-1:0]      phy_txeq_ctrl_o,      
   output wire [(PHY_LANE*4)-1:0]      phy_txeq_preset_o,       
   output wire [(PHY_LANE*6)-1:0]      phy_txeq_coeff_o,    

   input  wire [ 5:0]                  phy_txeq_fs_i,           
   input  wire [ 5:0]                  phy_txeq_lf_i,           
   input  wire [(PHY_LANE*18)-1:0]     phy_txeq_new_coeff_i,        
   input  wire [PHY_LANE-1:0]          phy_txeq_done_i,         

   output wire [ 5:0]                  phy_txeq_fs_o,           
   output wire [ 5:0]                  phy_txeq_lf_o,           
   output wire [(PHY_LANE*18)-1:0]     phy_txeq_new_coeff_o,        
   output wire [PHY_LANE-1:0]          phy_txeq_done_o,         

   // RX Equalization (Gen3/4)
   input  wire [(PHY_LANE*2)-1:0]      phy_rxeq_ctrl_i,     
   input  wire [(PHY_LANE*4)-1:0]      phy_rxeq_txpreset_i,   

   output wire [(PHY_LANE*2)-1:0]      phy_rxeq_ctrl_o,     
   output wire [(PHY_LANE*4)-1:0]      phy_rxeq_txpreset_o,      

   input  wire [PHY_LANE-1:0]          phy_rxeq_preset_sel_i,    
   input  wire [(PHY_LANE*18)-1:0]     phy_rxeq_new_txcoeff_i,   
   input  wire [PHY_LANE-1:0]          phy_rxeq_adapt_done_i,     
   input  wire [PHY_LANE-1:0]          phy_rxeq_done_i,

   output wire [PHY_LANE-1:0]          phy_rxeq_preset_sel_o,    
   output wire [(PHY_LANE*18)-1:0]     phy_rxeq_new_txcoeff_o,   
   output wire [PHY_LANE-1:0]          phy_rxeq_adapt_done_o,     
   output wire [PHY_LANE-1:0]          phy_rxeq_done_o,

   // Assist Signals
   input  wire                         as_mac_in_detect_i,
   input  wire                         as_cdr_hold_req_i,

   output wire                         as_mac_in_detect_o,
   output wire                         as_cdr_hold_req_o
   );

   genvar         lane;

generate
   for (lane = 0; lane < PHY_LANE; lane = lane + 1) begin: per_lane_ff_chain
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 64, 64'd0, phy_txdata_chain, phy_pclk, phy_rst, phy_txdata_o[(lane* 64)+:64], phy_txdata_i[(lane* 64)+:64])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 2, 2'd0, phy_txdatak_chain, phy_pclk, phy_rst, phy_txdatak_o[(lane* 2)+:2], phy_txdatak_i[(lane* 2)+:2])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd0, phy_txdata_valid_chain, phy_pclk, phy_rst, phy_txdata_valid_o[lane], phy_txdata_valid_i[lane])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd0, phy_txstart_block_chain, phy_pclk, phy_rst, phy_txstart_block_o[lane], phy_txstart_block_i[lane])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 2, 2'd0, phy_txsync_header_chain, phy_pclk, phy_rst, phy_txsync_header_o[(lane* 2)+:2], phy_txsync_header_i[(lane* 2)+:2])

      `FF_CHAIN_MODEL(PIPELINE_STAGES, 64, 64'd0, phy_rxdata_chain, phy_pclk, phy_rst, phy_rxdata_o[(lane* 64)+:64], phy_rxdata_i[(lane* 64)+:64])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 2, 2'd0, phy_rxdatak_chain, phy_pclk, phy_rst, phy_rxdatak_o[(lane* 2)+:2], phy_rxdatak_i[(lane* 2)+:2])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd0, phy_rxdata_valid_chain, phy_pclk, phy_rst, phy_rxdata_valid_o[lane], phy_rxdata_valid_i[lane])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 2, 2'd0, phy_rxstart_block_chain, phy_pclk, phy_rst, phy_rxstart_block_o[(lane* 2)+:2], phy_rxstart_block_i[(lane* 2)+:2])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 2, 2'd0, phy_rxsync_header_chain, phy_pclk, phy_rst, phy_rxsync_header_o[(lane* 2)+:2], phy_rxsync_header_i[(lane* 2)+:2])

      `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd1, phy_txelecidle_chain, phy_pclk, phy_rst, phy_txelecidle_o[lane], phy_txelecidle_i[lane])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd0, phy_txcompliance_chain, phy_pclk, phy_rst, phy_txcompliance_o[lane], phy_txcompliance_i[lane])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd0, phy_rxpolarity_chain, phy_pclk, phy_rst, phy_rxpolarity_o[lane], phy_rxpolarity_i[lane])

      `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd0, phy_rxvalid_chain, phy_pclk, phy_rst, phy_rxvalid_o[lane], phy_rxvalid_i[lane])
      `AS_FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd1, phy_phystatus_chain, phy_pclk, phy_rst, phy_phystatus_o[lane], phy_phystatus_i[lane])
      `AS_FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd1, phy_rxelecidle_chain, phy_pclk, phy_rst, phy_rxelecidle_o[lane], phy_rxelecidle_i[lane])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 3, 3'd0, phy_rxstatus_chain, phy_pclk, phy_rst, phy_rxstatus_o[(lane* 3)+:3], phy_rxstatus_i[(lane* 3)+:3])

      `FF_CHAIN_MODEL(PIPELINE_STAGES, 2, 2'd0, phy_txeq_ctrl_chain, phy_pclk, phy_rst, phy_txeq_ctrl_o[(lane* 2)+:2], phy_txeq_ctrl_i[(lane* 2)+:2])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 4, 6'd0, phy_txeq_preset_chain, phy_pclk, phy_rst, phy_txeq_preset_o[(lane* 4)+:4], phy_txeq_preset_i[(lane* 4)+:4])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 6, 6'd0, phy_txeq_coeff_chain, phy_pclk, phy_rst, phy_txeq_coeff_o[(lane* 6)+:6], phy_txeq_coeff_i[(lane* 6)+:6])

      `FF_CHAIN_MODEL(PIPELINE_STAGES,18,18'd0, phy_txeq_new_coeff_chain, phy_pclk, phy_rst, phy_txeq_new_coeff_o[(lane* 18)+:18], phy_txeq_new_coeff_i[(lane* 18)+:18])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd0, phy_txeq_done_chain, phy_pclk, phy_rst, phy_txeq_done_o[lane], phy_txeq_done_i[lane])

      `FF_CHAIN_MODEL(PIPELINE_STAGES, 2, 2'd0, phy_rxeq_ctrl_chain, phy_pclk, phy_rst, phy_rxeq_ctrl_o[(lane* 2)+:2], phy_rxeq_ctrl_i[(lane* 2)+:2])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 4, 6'd0, phy_rxeq_txpreset_chain, phy_pclk, phy_rst, phy_rxeq_txpreset_o[(lane* 4)+:4], phy_rxeq_txpreset_i[(lane* 4)+:4])

      `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd0, phy_rxeq_preset_sel_chain, phy_pclk, phy_rst, phy_rxeq_preset_sel_o[lane], phy_rxeq_preset_sel_i[lane])
      `FF_CHAIN_MODEL(PIPELINE_STAGES,18,18'd0, phy_rxeq_new_txcoeff_chain, phy_pclk, phy_rst, phy_rxeq_new_txcoeff_o[(lane* 18)+:18], phy_rxeq_new_txcoeff_i[(lane* 18)+:18])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd0, phy_rxeq_adapt_done_chain, phy_pclk, phy_rst, phy_rxeq_adapt_done_o[lane], phy_rxeq_adapt_done_i[lane])
      `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd0, phy_rxeq_done_chain, phy_pclk, phy_rst, phy_rxeq_done_o[lane], phy_rxeq_done_i[lane])
   end
endgenerate

   `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd0, phy_txdetectrx_chain, phy_pclk, phy_rst, phy_txdetectrx_o, phy_txdetectrx_i)
   `FF_CHAIN_MODEL(PIPELINE_STAGES, 2, 2'd2, phy_powerdown_chain, phy_pclk, phy_rst, phy_powerdown_o, phy_powerdown_i)
   `FF_CHAIN_MODEL(PIPELINE_STAGES, 2, 2'd0, phy_rate_chain, phy_pclk, phy_rst, phy_rate_o, phy_rate_i)
   `FF_CHAIN_MODEL(PIPELINE_STAGES, 3, 3'd0, phy_txmargin_chain, phy_pclk, phy_rst, phy_txmargin_o, phy_txmargin_i)
   `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd0, phy_txswing_chain, phy_pclk, phy_rst, phy_txswing_o, phy_txswing_i)
   `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd1, phy_txdeemph_chain, phy_pclk, phy_rst, phy_txdeemph_o, phy_txdeemph_i)
   `FF_CHAIN_MODEL(PIPELINE_STAGES, 6, 6'd0, phy_txeq_fs_chain, phy_pclk, phy_rst, phy_txeq_fs_o, phy_txeq_fs_i) 
   `FF_CHAIN_MODEL(PIPELINE_STAGES, 6, 6'd0, phy_txeq_lf_chain, phy_pclk, phy_rst, phy_txeq_lf_o, phy_txeq_lf_i)
   `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd1, as_mac_in_detect_chain, phy_pclk, phy_rst, as_mac_in_detect_o, as_mac_in_detect_i)
   `FF_CHAIN_MODEL(PIPELINE_STAGES, 1, 1'd0, as_cdr_hold_req_chain, phy_pclk, phy_rst, as_cdr_hold_req_o, as_cdr_hold_req_i)

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_pl_eq.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_pl_eq #(
    parameter             TCQ = 100
   ,parameter             IMPL_TARGET = "SOFT"
   ,parameter             PL_UPSTREAM_FACING="TRUE"
  ) (
   
    input  wire           clk_i
   ,input  wire           reset_i
   ,input  wire           link_down_reset_i

   ,input  wire [5:0]     cfg_ltssm_state_i
   ,input  wire           pl_redo_eq_i
   ,input  wire           pl_redo_eq_speed_i
   ,output reg            pl_eq_mismatch_o
   ,output reg            pl_redo_eq_pending_o
   
   ,output wire           pl_gen34_redo_equalization_o
   ,output wire           pl_gen34_redo_eq_speed_o
   ,input  wire           pl_gen34_eq_mismatch_i
   );

   reg                    pl_eq_mismatch_w;
   reg                    pl_redo_eq_pending_w;

   generate  
  
     if (PL_UPSTREAM_FACING == "TRUE") begin 

       always @(*) begin

         pl_eq_mismatch_w = pl_eq_mismatch_o;
         pl_redo_eq_pending_w = pl_redo_eq_pending_o;
    
         if (!pl_eq_mismatch_o && (cfg_ltssm_state_i[5:0] == 6'h0B) && pl_gen34_eq_mismatch_i) begin
    
           pl_eq_mismatch_w = 1'b1;
    
         end else if (!pl_redo_eq_pending_o && (cfg_ltssm_state_i[5:0] == 6'h0D) && pl_gen34_eq_mismatch_i) begin
    
           pl_redo_eq_pending_w = 1'b1;
      
         end else if (pl_redo_eq_pending_o && pl_redo_eq_i) begin
    
           pl_redo_eq_pending_w = 1'b0;
    
         end
    
       end

     end else begin // PL_UPSTREAM_FACING == FALSE
 
       always @(*) begin

         pl_eq_mismatch_w = pl_gen34_eq_mismatch_i;
         pl_redo_eq_pending_w = 1'b0;

       end

     end

   endgenerate
   
   always @(posedge clk_i) begin

     if (reset_i) begin

       pl_eq_mismatch_o <= #(TCQ) 1'b0;
       pl_redo_eq_pending_o <= #(TCQ) 1'b0;

     end else if (link_down_reset_i) begin   

       pl_eq_mismatch_o <= #(TCQ) 1'b0;
       pl_redo_eq_pending_o <= #(TCQ) 1'b0;

     end else begin
     
       pl_eq_mismatch_o <= #(TCQ) pl_eq_mismatch_w;
       pl_redo_eq_pending_o <= #(TCQ) pl_redo_eq_pending_w;

     end

   end

   assign pl_gen34_redo_equalization_o = pl_redo_eq_i;
   assign pl_gen34_redo_eq_speed_o = pl_redo_eq_speed_i;

endmodule // pcie_4_0_pl_eq
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_seqnum_fifo.v
// Version    : 1.1 
//-----------------------------------------------------------------------------

`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_seqnum_fifo #(

  // Parameters

  parameter            TCQ                               = 1,
  parameter 		       RAM_WIDTH                         = 6,
  parameter 		       RAM_DEPTH                         = 4,
  parameter 		       ADDR_WIDTH                        = 2,
  parameter 		       FIFO_FULL_HIGH_THRESHOLD          = 3'd4,
  parameter 		       FIFO_FULL_LOW_THRESHOLD           = 3'd1,

  parameter 		       IN_FSM_SIZE                       = 2,
  parameter 		       IN_FSM_IDLE                       = 2'b01,
  parameter 		       IN_FSM_CHANGE                     = 2'b10,
  parameter            NO_UPDATE_PREV_DATA_ON_FIFO_FULL  = 1'b0
  )
  (
  input 	                    core_reset_n_i,
  input                       core_clk_i,

  input                       user_reset_n_i,
  input                       user_clk_i,

  input  [(RAM_WIDTH-1):0]    data_i, 
  output [(RAM_WIDTH-1):0]    data_o

  );  


  // Local Registers

  reg [RAM_WIDTH-1:0] 	       reg_ram[RAM_DEPTH-1:0];

  integer                      index;
  reg [ADDR_WIDTH:0] 	       write_addr;
  reg [ADDR_WIDTH:0] 	       write_addr_read_clk;
  reg [ADDR_WIDTH:0] 	       read_addr;
  reg [ADDR_WIDTH:0] 	       read_addr_wrclk;
  reg 			       fifo_full;

  reg [(IN_FSM_SIZE-1):0]      reg_in_fsm_state /* synthesis syn_state_machine=1 */;
  reg [(IN_FSM_SIZE-1):0]      reg_in_fsm_next_state;

  reg [(RAM_WIDTH-1):0]        reg_prev_data;
  reg [(RAM_WIDTH-1):0]        reg_out_data;

  reg [(RAM_WIDTH-1):0]        data_int;

  // Local wires

  wire [ADDR_WIDTH:0] 	       write_addr_next;
  wire [ADDR_WIDTH:0] 	       read_addr_next;
  wire [ADDR_WIDTH:0] 	       read_side_occupancy;
  wire [ADDR_WIDTH:0] 	       write_side_occupancy;
  wire 			       read_data_valid;
  wire 			       fifo_empty;
  wire 			       write_enable;
  wire [RAM_WIDTH-1:0] 	       ram_write_data;
  wire [RAM_WIDTH-1:0] 	       ram_read_data;

  wire [(RAM_WIDTH-1):0]       prev_data_w;
 
  wire [(IN_FSM_SIZE-1):0]     in_fsm_state_w;

  //  Capture data_i
  always @(posedge core_clk_i or negedge core_reset_n_i)
    if (~core_reset_n_i)
      data_int <= #(TCQ) {RAM_WIDTH{1'b0}};
    else 
      data_int <= #(TCQ) data_i;

  // Capture LTSSM state on change
  always @(posedge core_clk_i or negedge core_reset_n_i)
    if (~core_reset_n_i)
      reg_prev_data <= #(TCQ) {RAM_WIDTH{1'b0}};
    else if (((data_int != prev_data_w) || (in_fsm_state_w == IN_FSM_CHANGE) ) & 
	     (~NO_UPDATE_PREV_DATA_ON_FIFO_FULL | (~fifo_full & NO_UPDATE_PREV_DATA_ON_FIFO_FULL)))
      reg_prev_data <= #(TCQ) data_int;
  
  // FSM Looks for change in the LTSSM state

  always @(posedge core_clk_i or negedge core_reset_n_i)
    if (~core_reset_n_i)
      reg_in_fsm_state <= #(TCQ) IN_FSM_IDLE;
    else
      reg_in_fsm_state <= #(TCQ) reg_in_fsm_next_state;

  // FSM Next State Logic

  always @( * )
    case (in_fsm_state_w)
      IN_FSM_IDLE :
        if (data_int != reg_prev_data)
          reg_in_fsm_next_state = IN_FSM_CHANGE;
        else
          reg_in_fsm_next_state = IN_FSM_IDLE;
      IN_FSM_CHANGE : 
        reg_in_fsm_next_state = IN_FSM_IDLE;
      default : 
        reg_in_fsm_next_state = IN_FSM_IDLE;
    endcase   

  // FIFO Write Side Processes

  assign  ram_write_data = data_int;
  //assign  write_enable = (data_int != prev_data_w) || (in_fsm_state_w == IN_FSM_CHANGE);
  assign  write_enable = (data_int[6]);
  assign  write_addr_next = write_addr + {{ADDR_WIDTH{1'b0}}, 1'b1};

  always @(posedge core_clk_i or negedge core_reset_n_i)
    if (~core_reset_n_i)
      write_addr <= {ADDR_WIDTH+1{1'b0}};
    else if (write_enable & ~fifo_full)
      write_addr <= write_addr_next;

  // Write into RAM 
  always @(posedge core_clk_i or negedge core_reset_n_i)
    if (~core_reset_n_i)
      begin
	for (index=0; index < RAM_DEPTH; index=index+1)
	  reg_ram[index] <= {RAM_WIDTH{1'b0}};
      end
    else if (write_enable)
      reg_ram[write_addr[ADDR_WIDTH-1:0]] <= ram_write_data;

  // FIFO Read Side Processes

  assign      read_addr_next = read_addr +  {{ADDR_WIDTH-1{1'b0}}, 1'b1};

  always @(posedge user_clk_i or negedge user_reset_n_i)
    if (~user_reset_n_i)
      read_addr <= {ADDR_WIDTH+1{1'b0}};
    else if (read_data_valid)
      read_addr <= read_addr_next;

  // Convert write pointer to the read clk domain
  always @(posedge user_clk_i or negedge user_reset_n_i)
    if (~user_reset_n_i)
      write_addr_read_clk <= {ADDR_WIDTH+1{1'b0}};
    else
      write_addr_read_clk <= write_addr;
  
  // Maintain read-side occupancy
  assign read_side_occupancy = (write_addr_read_clk - read_addr);
  assign fifo_empty = (read_side_occupancy == {ADDR_WIDTH+1{1'b0}});
  assign read_data_valid = ~fifo_empty;
  assign ram_read_data = reg_ram[read_addr[ADDR_WIDTH-1:0]];

  /* convert read pointer to write clock domain */
  always @(posedge core_clk_i or negedge core_reset_n_i)
    if (~core_reset_n_i)
      read_addr_wrclk <= {ADDR_WIDTH+1{1'b0}};
    else
      read_addr_wrclk <= read_addr;

  assign write_side_occupancy = write_addr - read_addr_wrclk;

  // Generate FIFO full condition
  always @(posedge core_clk_i or negedge core_reset_n_i)
    if (~core_reset_n_i)
      fifo_full <= 1'b0;
    else
      if (write_side_occupancy[ADDR_WIDTH] ||
	  (write_side_occupancy[ADDR_WIDTH-1:0] == FIFO_FULL_HIGH_THRESHOLD))
	fifo_full <= 1'b1;
      else
	// Clear when FIFO occupancy goes below low threshold
	if (~write_side_occupancy[ADDR_WIDTH] &&
	    (write_side_occupancy[ADDR_WIDTH-1:0] <= FIFO_FULL_LOW_THRESHOLD))
	  fifo_full <= 1'b0;

  // Latch Last
  always @(posedge user_clk_i or negedge user_reset_n_i)
    if (~user_reset_n_i)
      reg_out_data <= #(TCQ) {RAM_WIDTH{1'b0}};
    else
      if (read_data_valid)
        reg_out_data <= #(TCQ) ram_read_data;
      else
	reg_out_data <= #(TCQ) 'h0;

  // Assignments

  assign in_fsm_state_w = reg_in_fsm_state;
  assign data_o = reg_out_data;
  assign prev_data_w = reg_prev_data; 
  
endmodule // pcie3_ccm_fifo
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_vf_decode.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_vf_decode #(

  parameter           TCQ = 100
 ,parameter           NUM_VFS = 252
 ,parameter [1:0]     TL_PF_ENABLE_REG=2'h0
 ,parameter [15:0]    PF0_SRIOV_CAP_TOTAL_VF=16'h0
 ,parameter [15:0]    PF1_SRIOV_CAP_TOTAL_VF=16'h0
 ,parameter [15:0]    PF2_SRIOV_CAP_TOTAL_VF=16'h0
 ,parameter [15:0]    PF3_SRIOV_CAP_TOTAL_VF=16'h0
 ,parameter [15:0]    PF0_SRIOV_FIRST_VF_OFFSET=16'h0
 ,parameter [15:0]    PF1_SRIOV_FIRST_VF_OFFSET=16'h0
 ,parameter [15:0]    PF2_SRIOV_FIRST_VF_OFFSET=16'h0
 ,parameter [15:0]    PF3_SRIOV_FIRST_VF_OFFSET=16'h0
 ,parameter [3:0]     SRIOV_CAP_ENABLE=4'h0
 ,parameter           ARI_CAP_ENABLE="FALSE"


  ) (

  input wire          clk_i
 ,input wire          reset_i
 ,input wire          link_down_i
 ,input wire          cfg_ext_write_received_i
 ,input wire [9:0]    cfg_ext_register_number_i
 ,input wire [7:0]    cfg_ext_function_number_i
 ,input wire [31:0]   cfg_ext_write_data_i
 ,input wire [3:0]    cfg_ext_write_byte_enable_i
 ,input wire [3:0]    cfg_flr_in_process_i

 ,output reg [NUM_VFS-1:0]   cfg_vf_flr_in_process_o
 ,output reg [2*NUM_VFS-1:0] cfg_vf_status_o          // Bit 0: Memory Space Enable; Bit 1: Bus Master Enable
 ,output reg [3*NUM_VFS-1:0] cfg_vf_power_state_o     // 000b - D0-Uninitialized; 001b - D0-Active; 010b - D1; 100b - D3hot
 ,output reg [NUM_VFS-1:0]   cfg_vf_tph_requester_enable_o
 ,output reg [3*NUM_VFS-1:0] cfg_vf_tph_st_mode_o     
 ,output reg [NUM_VFS-1:0]   cfg_interrupt_msix_vf_enable_o
 ,output reg [NUM_VFS-1:0]   cfg_interrupt_msix_vf_mask_o

  );

  localparam [9:0]   REG_DEV_CTRL=10'h1E;
  localparam         REG_DEV_CTRL__FLR_SIZE=1;
  localparam         REG_DEV_CTRL__FLR=15;

  localparam [9:0]   REG_PCI_CMD=10'h1;
  localparam         REG_PCI_CMD__BME_SIZE=1;  
  localparam         REG_PCI_CMD__BME=2;
  localparam         REG_PCI_CMD__MSE_SIZE=1;  
  localparam         REG_PCI_CMD__MSE=1;  

  localparam [9:0]   REG_PM_CSR=10'h11;
  localparam         REG_PM_CSR__PS_SIZE=2;
  localparam         REG_PM_CSR__PS=0;

  localparam [9:0]   REG_TPH_CR=10'h8A;
  localparam         REG_TPH_CR__RQE_SIZE=1;  
  localparam         REG_TPH_CR__RQE=8;  
  localparam         REG_TPH_CR__STMS_SIZE=3;
  localparam         REG_TPH_CR__STMS=0;

  localparam [9:0]   REG_MSIX_CR=10'h18;
  localparam         REG_MSIX_CR__EN_SIZE=1;  
  localparam         REG_MSIX_CR__EN=31;  
  localparam         REG_MSIX_CR__MSK_SIZE=1;
  localparam         REG_MSIX_CR__MSK=30;
  localparam         PF_VF_MAP_WIDTH=256;

  reg                 cfg_ext_write_received;
  reg [9:0]           cfg_ext_register_number;
  reg [7:0]           cfg_ext_function_number;
  reg [31:0]          cfg_ext_write_data;
  reg [3:0]           cfg_ext_write_byte_enable;

  reg [NUM_VFS-1:0]   cfg_vf_flr_in_process_w;
  reg [2*NUM_VFS-1:0] cfg_vf_status_w;
  reg [3*NUM_VFS-1:0] cfg_vf_power_state_w;
  reg [NUM_VFS-1:0]   cfg_vf_tph_requester_enable_w;
  reg [3*NUM_VFS-1:0] cfg_vf_tph_st_mode_w;
  reg [NUM_VFS-1:0]   cfg_interrupt_msix_vf_enable_w;
  reg [NUM_VFS-1:0]   cfg_interrupt_msix_vf_mask_w;
  reg [NUM_VFS-1:0]   cfg_interrupt_msix_vf_flr_msk_w;
  reg [NUM_VFS-1:0]   reg_cfg_interrupt_msix_vf_flr_msk;

  wire [NUM_VFS-1:0]  cfg_vf_active_w;
  reg [NUM_VFS-1:0]   reg_cfg_vf_active;
  reg [NUM_VFS-1:0]   cfg_vf_active;

  wire [7:0]          cfg_ext_function_number_w;
  wire [7:0]          cfg_ext_function_number_w_2_b0;
  wire [7:0]          cfg_ext_function_number_w_2_b1;
  wire [7:0]          cfg_ext_function_number_w_3_b0;
  wire [7:0]          cfg_ext_function_number_w_3_b1;
  wire [7:0]          cfg_ext_function_number_w_3_b2;
  wire [3:0]          pf_mapenable;
  wire                pf_as_vf;
  wire [2:0]          pf_as_vf_mapd;

  // Only use attributes in these static assignments for PF_VF_MAP
  wire [(PF_VF_MAP_WIDTH-1):0] pf0_vf_size;
  wire [(PF_VF_MAP_WIDTH-1):0] pf1_vf_size;
  wire [(PF_VF_MAP_WIDTH-1):0] pf2_vf_size;
  wire [(PF_VF_MAP_WIDTH-1):0] pf3_vf_size;
  wire [(PF_VF_MAP_WIDTH-1):0] pf0_vf_mapd;
  wire [(PF_VF_MAP_WIDTH-1):0] pf1_vf_mapd;
  wire [(PF_VF_MAP_WIDTH-1):0] pf2_vf_mapd;
  wire [(PF_VF_MAP_WIDTH-1):0] pf3_vf_mapd;

  wire [(PF_VF_MAP_WIDTH-1):0] pf0_vf_map_w;
  wire [(PF_VF_MAP_WIDTH-1):0] pf1_vf_map_w;
  wire [(PF_VF_MAP_WIDTH-1):0] pf2_vf_map_w;
  wire [(PF_VF_MAP_WIDTH-1):0] pf3_vf_map_w;

  integer                      i;

  always @(posedge clk_i) begin
  
    if (reset_i) begin

      cfg_ext_write_received <= #(TCQ) 1'b0;
      cfg_ext_register_number <= #(TCQ) 10'b0;
      cfg_ext_function_number <= #(TCQ) 8'b0;
      cfg_ext_write_data <= #(TCQ) 32'b0;
      cfg_ext_write_byte_enable <= #(TCQ) 4'b0;

      cfg_vf_flr_in_process_o <= #(TCQ) {NUM_VFS{1'b0}};
      cfg_vf_status_o <= #(TCQ) {2*NUM_VFS{1'b0}};
      cfg_vf_power_state_o <= #(TCQ) {3*NUM_VFS{1'b0}};
      cfg_vf_tph_requester_enable_o <= #(TCQ) {2*NUM_VFS{1'b0}};
      cfg_vf_tph_st_mode_o <= #(TCQ) {3*NUM_VFS{1'b0}};
      cfg_interrupt_msix_vf_enable_o <= #(TCQ) {NUM_VFS{1'b0}};
      cfg_interrupt_msix_vf_mask_o <= #(TCQ) {NUM_VFS{1'b0}};

      reg_cfg_vf_active <= #(TCQ) {NUM_VFS{1'b0}};
      reg_cfg_interrupt_msix_vf_flr_msk <= #(TCQ) {NUM_VFS{1'b1}};   

    end else if (link_down_i) begin

      cfg_ext_write_received <= #(TCQ) 1'b0;
      cfg_ext_register_number <= #(TCQ) 10'b0;
      cfg_ext_function_number <= #(TCQ) 8'b0;
      cfg_ext_write_data <= #(TCQ) 32'b0;
      cfg_ext_write_byte_enable <= #(TCQ) 4'b0;

      cfg_vf_flr_in_process_o <= #(TCQ) {NUM_VFS{1'b0}};
      cfg_vf_status_o <= #(TCQ) {2*NUM_VFS{1'b0}};
      cfg_vf_power_state_o <= #(TCQ) {3*NUM_VFS{1'b0}};
      cfg_vf_tph_requester_enable_o <= #(TCQ) {2*NUM_VFS{1'b0}};
      cfg_vf_tph_st_mode_o <= #(TCQ) {3*NUM_VFS{1'b0}};
      cfg_interrupt_msix_vf_enable_o <= #(TCQ) {NUM_VFS{1'b0}};
      cfg_interrupt_msix_vf_mask_o <= #(TCQ) {NUM_VFS{1'b0}};

      reg_cfg_vf_active <= #(TCQ) {NUM_VFS{1'b0}};
      reg_cfg_interrupt_msix_vf_flr_msk <= #(TCQ) {NUM_VFS{1'b1}};   

    end else begin

      cfg_ext_write_received <= #(TCQ) cfg_ext_write_received_i;
      cfg_ext_register_number <= #(TCQ) cfg_ext_register_number_i;
      cfg_ext_function_number <= #(TCQ) cfg_ext_function_number_i; 
      cfg_ext_write_data <= #(TCQ) cfg_ext_write_data_i;
      cfg_ext_write_byte_enable <= #(TCQ) cfg_ext_write_byte_enable_i;

      cfg_vf_flr_in_process_o <= #(TCQ) cfg_vf_flr_in_process_w;
      cfg_vf_status_o <= #(TCQ) cfg_vf_status_w;
      cfg_vf_power_state_o <= #(TCQ) cfg_vf_power_state_w;
      cfg_vf_tph_requester_enable_o <= #(TCQ) cfg_vf_tph_requester_enable_w;
      cfg_vf_tph_st_mode_o <= #(TCQ) cfg_vf_tph_st_mode_w;
      cfg_interrupt_msix_vf_enable_o <= #(TCQ) cfg_interrupt_msix_vf_enable_w & cfg_interrupt_msix_vf_flr_msk_w;
      cfg_interrupt_msix_vf_mask_o <= #(TCQ) cfg_interrupt_msix_vf_mask_w & cfg_interrupt_msix_vf_flr_msk_w;

      reg_cfg_vf_active <= #(TCQ) cfg_vf_active_w;
      reg_cfg_interrupt_msix_vf_flr_msk <= #(TCQ) cfg_interrupt_msix_vf_flr_msk_w;

    end

  end

  /*
  *  1)
  *  if any of the PF sees a FLR (cfg_flr_in_process_i bits set to 1b),
  *  then, corresponding VF bits in cfg_interrupt_msix_vf_enable_o and
  *  cfg_interrupt_msix_vf_mask_o must be reset.
  *  2)
  *  if any of the VF sees a FLR (cfg_vf_flr_in_process_w bits set to 1b),
  *  then, corresponding VF bits in cfg_interrupt_msix_vf_enable_o and
  *  cfg_interrupt_msix_vf_mask_o must be reset.
  */

  always @ (*) begin

    for (i = 0; i < 252; i = i + 1) begin

      if (cfg_flr_in_process_i[0] & pf0_vf_map_w[i+4])
        cfg_interrupt_msix_vf_flr_msk_w[i] = 1'b0;
      else if (!cfg_flr_in_process_i[0] & pf0_vf_map_w[i+4])
        cfg_interrupt_msix_vf_flr_msk_w[i] = 1'b1;
      else
	cfg_interrupt_msix_vf_flr_msk_w[i] = reg_cfg_interrupt_msix_vf_flr_msk[i];

    end

    for (i = 0; i < 252; i = i + 1) begin

      if (cfg_flr_in_process_i[1] & pf1_vf_map_w[i+4])
        cfg_interrupt_msix_vf_flr_msk_w[i] = 1'b0; 
      else if (!cfg_flr_in_process_i[1] & pf1_vf_map_w[i+4])
        cfg_interrupt_msix_vf_flr_msk_w[i] = 1'b1; 
      else
	cfg_interrupt_msix_vf_flr_msk_w[i] = reg_cfg_interrupt_msix_vf_flr_msk[i];

    end

    for (i = 0; i < 252; i = i + 1) begin

      if (cfg_flr_in_process_i[2] & pf2_vf_map_w[i+4])
        cfg_interrupt_msix_vf_flr_msk_w[i] = 1'b0; 
      else if (!cfg_flr_in_process_i[2] & pf2_vf_map_w[i+4])
        cfg_interrupt_msix_vf_flr_msk_w[i] = 1'b1; 
      else
	cfg_interrupt_msix_vf_flr_msk_w[i] = reg_cfg_interrupt_msix_vf_flr_msk[i];

    end

    for (i = 0; i < 252; i = i + 1) begin

      if (cfg_flr_in_process_i[3] & pf3_vf_map_w[i+4])
        cfg_interrupt_msix_vf_flr_msk_w[i] = 1'b0; 
      else if (!cfg_flr_in_process_i[3] & pf3_vf_map_w[i+4])
        cfg_interrupt_msix_vf_flr_msk_w[i] = 1'b1; 
      else
	cfg_interrupt_msix_vf_flr_msk_w[i] = reg_cfg_interrupt_msix_vf_flr_msk[i];

    end

    for (i = 0; i < 252; i = i + 1) begin

      if (cfg_vf_flr_in_process_w[i])
        cfg_interrupt_msix_vf_flr_msk_w[i] = 1'b0;
      else
        cfg_interrupt_msix_vf_flr_msk_w[i] = 1'b1;

    end

  end

  always @(*) begin

    cfg_vf_flr_in_process_w = cfg_vf_flr_in_process_o;
    cfg_vf_status_w = cfg_vf_status_o;
    cfg_vf_power_state_w = cfg_vf_power_state_o;
    cfg_vf_tph_requester_enable_w = cfg_vf_tph_requester_enable_o;
    cfg_vf_tph_st_mode_w = cfg_vf_tph_st_mode_o;
    cfg_interrupt_msix_vf_enable_w = cfg_interrupt_msix_vf_enable_o; 
    cfg_interrupt_msix_vf_mask_w = cfg_interrupt_msix_vf_mask_o;
    cfg_vf_active = cfg_vf_active_w;

    if (cfg_ext_write_received && (cfg_ext_function_number > 3)) begin

      if (cfg_ext_register_number == REG_DEV_CTRL) begin

        if (cfg_ext_write_byte_enable[1])
          cfg_vf_flr_in_process_w[cfg_ext_function_number_w] = cfg_ext_write_data[REG_DEV_CTRL__FLR];

      end else if (cfg_ext_register_number == REG_PCI_CMD) begin

        if (cfg_ext_write_byte_enable[0]) begin

          cfg_vf_status_w[cfg_ext_function_number_w_2_b0] = cfg_ext_write_data[REG_PCI_CMD__MSE]; 
          cfg_vf_status_w[cfg_ext_function_number_w_2_b1] = cfg_ext_write_data[REG_PCI_CMD__BME]; 
          cfg_vf_active[cfg_ext_function_number_w] = cfg_ext_write_data[REG_PCI_CMD__BME] | cfg_ext_write_data[REG_PCI_CMD__MSE];
          // if Function in D0-Uninit then transtion to D0-Active
          if ((!cfg_vf_power_state_w[cfg_ext_function_number_w_3_b0]) &&
              (!cfg_vf_power_state_w[cfg_ext_function_number_w_3_b1]) &&
              (!cfg_vf_power_state_w[cfg_ext_function_number_w_3_b2]))
            cfg_vf_power_state_w[cfg_ext_function_number_w_3_b0] = cfg_vf_active_w[cfg_ext_function_number_w];

        end

      end else if (cfg_ext_register_number == REG_PM_CSR) begin

        if (cfg_ext_write_byte_enable[0]) begin

          cfg_vf_power_state_w[cfg_ext_function_number_w_3_b0] = cfg_vf_active[cfg_ext_function_number_w] && 
					                           (!cfg_ext_write_data[REG_PM_CSR__PS] || 
					                            !cfg_ext_write_data[REG_PM_CSR__PS+REG_PM_CSR__PS_SIZE-1]);
          cfg_vf_power_state_w[cfg_ext_function_number_w_3_b1] = (cfg_ext_write_data[REG_PM_CSR__PS] && 
		                                                  !cfg_ext_write_data[REG_PM_CSR__PS+REG_PM_CSR__PS_SIZE-1]); 
          cfg_vf_power_state_w[cfg_ext_function_number_w_3_b2] = (cfg_ext_write_data[REG_PM_CSR__PS] && 
		                                                  cfg_ext_write_data[REG_PM_CSR__PS+REG_PM_CSR__PS_SIZE-1]); 

        end

      end else if (cfg_ext_register_number == REG_TPH_CR) begin

        if (cfg_ext_write_byte_enable[0]) begin

          cfg_vf_tph_st_mode_w[cfg_ext_function_number_w_3_b0] = cfg_ext_write_data[REG_TPH_CR__STMS];
          cfg_vf_tph_st_mode_w[cfg_ext_function_number_w_3_b1] = cfg_ext_write_data[REG_TPH_CR__STMS+1]; 
          cfg_vf_tph_st_mode_w[cfg_ext_function_number_w_3_b2] = cfg_ext_write_data[REG_TPH_CR__STMS+2]; 

        end

        if (cfg_ext_write_byte_enable[1])
          cfg_vf_tph_requester_enable_w[cfg_ext_function_number_w] = cfg_ext_write_data[REG_TPH_CR__RQE]; 

      end else if (cfg_ext_register_number == REG_MSIX_CR) begin

        if (cfg_ext_write_byte_enable[3]) begin
          cfg_interrupt_msix_vf_enable_w[cfg_ext_function_number_w] = cfg_ext_write_data[REG_MSIX_CR__EN];
          cfg_interrupt_msix_vf_mask_w[cfg_ext_function_number_w] = cfg_ext_write_data[REG_MSIX_CR__MSK];
        end

      end

    end

  end

  assign cfg_ext_function_number_w = cfg_ext_function_number - 4;
  assign cfg_ext_function_number_w_2_b0 = 2*(cfg_ext_function_number_w)+0;
  assign cfg_ext_function_number_w_2_b1 = 2*(cfg_ext_function_number_w)+1;
  assign cfg_ext_function_number_w_3_b0 = 3*(cfg_ext_function_number_w)+0;
  assign cfg_ext_function_number_w_3_b1 = 3*(cfg_ext_function_number_w)+1;
  assign cfg_ext_function_number_w_3_b2 = 3*(cfg_ext_function_number_w)+2;
  assign cfg_vf_active_w = reg_cfg_vf_active;

  // Decoded number of pfs
  assign pf_mapenable[0] = 1'b1;
  assign pf_mapenable[1] = (TL_PF_ENABLE_REG == 2'h1) | (TL_PF_ENABLE_REG == 2'h2) | (TL_PF_ENABLE_REG == 2'h3) ;
  assign pf_mapenable[2] = (TL_PF_ENABLE_REG == 2'h2) | (TL_PF_ENABLE_REG == 2'h3) ;
  assign pf_mapenable[3] = (TL_PF_ENABLE_REG == 2'h3) ;
  
  // These bit-widths are sized for max. 256 functions and single bus no.
  assign pf0_vf_size = {PF_VF_MAP_WIDTH{pf_mapenable[0]}} << PF0_SRIOV_CAP_TOTAL_VF[7:0];
  assign pf1_vf_size = {PF_VF_MAP_WIDTH{pf_mapenable[1]}} << PF1_SRIOV_CAP_TOTAL_VF[7:0];
  assign pf2_vf_size = {PF_VF_MAP_WIDTH{pf_mapenable[2]}} << PF2_SRIOV_CAP_TOTAL_VF[7:0];
  assign pf3_vf_size = {PF_VF_MAP_WIDTH{pf_mapenable[3]}} << PF3_SRIOV_CAP_TOTAL_VF[7:0];
  
  // Make sure to disable the VFs based on the individual PF enables
  assign pf0_vf_mapd = pf_mapenable[0] ? (~pf0_vf_size << (        PF0_SRIOV_FIRST_VF_OFFSET[7:0])) : 'b0;
  assign pf1_vf_mapd = pf_mapenable[1] ? (~pf1_vf_size << (8'h01 + PF1_SRIOV_FIRST_VF_OFFSET[7:0])) : 'b0;
  assign pf2_vf_mapd = pf_mapenable[2] ? (~pf2_vf_size << (8'h02 + PF2_SRIOV_FIRST_VF_OFFSET[7:0])) : 'b0;
  assign pf3_vf_mapd = pf_mapenable[3] ? (~pf3_vf_size << (8'h03 + PF3_SRIOV_FIRST_VF_OFFSET[7:0])) : 'b0;
  
  assign pf_as_vf = ((SRIOV_CAP_ENABLE[0] == 1'b1) && (ARI_CAP_ENABLE == "FALSE")) ;
  assign pf_as_vf_mapd = pf_as_vf ? pf0_vf_mapd[3:1] : 3'h0;
  
  assign pf0_vf_map_w = {pf0_vf_mapd[(PF_VF_MAP_WIDTH-1):4],{pf_as_vf_mapd,pf_mapenable[0]}};
  assign pf1_vf_map_w = {pf1_vf_mapd[(PF_VF_MAP_WIDTH-1):4],{2'h0,pf_mapenable[1],1'h0}};
  assign pf2_vf_map_w = {pf2_vf_mapd[(PF_VF_MAP_WIDTH-1):4],{1'h0,pf_mapenable[2],2'h0}};
  assign pf3_vf_map_w = {pf3_vf_mapd[(PF_VF_MAP_WIDTH-1):4],{pf_mapenable[3], 3'h0}};

endmodule



//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_bram.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_bram #(
  parameter           TCQ = 100
, parameter           AXISTEN_IF_MSIX_TO_RAM_PIPELINE="FALSE"
, parameter           AXISTEN_IF_MSIX_FROM_RAM_PIPELINE="FALSE"
, parameter           TPH_TO_RAM_PIPELINE="FALSE"
, parameter           TPH_FROM_RAM_PIPELINE="FALSE"
, parameter [1:0]     TL_COMPLETION_RAM_SIZE=2'b01
, parameter           TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE="FALSE"
, parameter           TL_RX_COMPLETION_TO_RAM_READ_PIPELINE="FALSE"
, parameter           TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE="FALSE"
, parameter           TL_RX_POSTED_TO_RAM_WRITE_PIPELINE="FALSE"
, parameter           TL_RX_POSTED_TO_RAM_READ_PIPELINE="FALSE"
, parameter           TL_RX_POSTED_FROM_RAM_READ_PIPELINE="FALSE"
, parameter           LL_REPLAY_TO_RAM_PIPELINE="FALSE"
, parameter           LL_REPLAY_FROM_RAM_PIPELINE="FALSE"
, parameter [1:0]     TL_PF_ENABLE_REG=2'h0
, parameter [3:0]     SRIOV_CAP_ENABLE=4'h0
, parameter [15:0]    PF0_SRIOV_CAP_TOTAL_VF=16'h0
, parameter [15:0]    PF1_SRIOV_CAP_TOTAL_VF=16'h0
, parameter [15:0]    PF2_SRIOV_CAP_TOTAL_VF=16'h0
, parameter [15:0]    PF3_SRIOV_CAP_TOTAL_VF=16'h0
, parameter           PF0_TPHR_CAP_ENABLE="FALSE"
, parameter           MSIX_CAP_TABLE_SIZE=11'h0
, parameter           MSIX_TABLE_RAM_ENABLE="FALSE"

  ) (
  input  wire         core_clk_i,
  input  wire         user_clk_i,
  input  wire         reset_i,

  input  wire   [8:0] mi_rep_addr_i,
  input  wire [255:0] mi_rep_wdata_i,
  input  wire         mi_rep_wen_i,
  output wire [255:0] mi_rep_rdata_o,
  input  wire         mi_rep_rden_i,

  output wire   [3:0] mi_rep_err_cor_o,
  output wire   [3:0] mi_rep_err_uncor_o,

  input  wire   [8:0] mi_req_waddr0_i,
  input  wire [143:0] mi_req_wdata0_i,
  input  wire         mi_req_wen0_i,
  input  wire   [8:0] mi_req_waddr1_i,
  input  wire [143:0] mi_req_wdata1_i,
  input  wire         mi_req_wen1_i,

  input  wire   [8:0] mi_req_raddr0_i,
  input  wire         mi_req_ren0_i,
  output wire [143:0] mi_req_rdata0_o,
  input  wire   [8:0] mi_req_raddr1_i,
  input  wire         mi_req_ren1_i,
  output wire [143:0] mi_req_rdata1_o,

  output wire   [5:0] mi_req_err_cor_o,
  output wire   [5:0] mi_req_err_uncor_o,

  input  wire   [8:0] mi_cpl_waddr0_i,
  input  wire [143:0] mi_cpl_wdata0_i,
  input  wire   [1:0] mi_cpl_wen0_i,
  input  wire   [8:0] mi_cpl_waddr1_i,
  input  wire [143:0] mi_cpl_wdata1_i,
  input  wire   [1:0] mi_cpl_wen1_i,

  input  wire   [8:0] mi_cpl_raddr0_i,
  input  wire   [1:0] mi_cpl_ren0_i,
  output wire [143:0] mi_cpl_rdata0_o,
  input  wire   [8:0] mi_cpl_raddr1_i,
  input  wire   [1:0] mi_cpl_ren1_i,
  output wire [143:0] mi_cpl_rdata1_o,

  output wire  [11:0] mi_cpl_err_cor_o,
  output wire  [11:0] mi_cpl_err_uncor_o,

  input  wire  [12:0] cfg_msix_waddr_i,
  input  wire  [31:0] cfg_msix_wdata_i,
  input  wire   [3:0] cfg_msix_wdip_i,
  input  wire   [3:0] cfg_msix_wen_i,
  output wire  [31:0] cfg_msix_rdata_o,
  output wire   [3:0] cfg_msix_rdop_o,
  input  wire         cfg_msix_ren_i,

  input  wire   [7:0] user_tph_stt_func_num_i,
  input  wire   [5:0] user_tph_stt_index_i,
  input  wire         user_tph_stt_rd_en_i,
  output wire   [7:0] user_tph_stt_rd_data_o,

  input  wire  [11:0] cfg_tph_waddr_i,
  input  wire  [31:0] cfg_tph_wdata_i,
  input  wire   [3:0] cfg_tph_wdip_i,
  input  wire   [3:0] cfg_tph_wen_i,
  output wire  [31:0] cfg_tph_rdata_o,
  output wire   [3:0] cfg_tph_rdop_o,
  input  wire         cfg_tph_ren_i

  );

  xp4_usp_smsw_bram_rep #(

    .TCQ (TCQ),
    .TO_RAM_PIPELINE(LL_REPLAY_TO_RAM_PIPELINE),
    .FROM_RAM_PIPELINE(LL_REPLAY_FROM_RAM_PIPELINE)

  )
  bram_repl_inst (

    .clk_i (core_clk_i),
    .reset_i (reset_i),

    .addr_i(mi_rep_addr_i[8:0]),
    .wdata_i(mi_rep_wdata_i[255:0]),
    .wen_i(mi_rep_wen_i),
    .rdata_o(mi_rep_rdata_o[255:0]),
    .ren_i(mi_rep_rden_i),
    .err_cor_o(mi_rep_err_cor_o[3:0]),
    .err_uncor_o(mi_rep_err_uncor_o[3:0])

  );

  xp4_usp_smsw_bram_16k #(

    .TCQ (TCQ),
    .TO_RAM_WRITE_PIPELINE(TL_RX_POSTED_TO_RAM_WRITE_PIPELINE),
    .TO_RAM_READ_PIPELINE(TL_RX_POSTED_TO_RAM_READ_PIPELINE),
    .FROM_RAM_READ_PIPELINE(TL_RX_POSTED_FROM_RAM_READ_PIPELINE)

  )
  bram_post_inst (

    .clk_i (core_clk_i),
    .reset_i (reset_i),

    .waddr0_i(mi_req_waddr0_i[8:0]),
    .wdata0_i(mi_req_wdata0_i[143:0]),
    .wen0_i(mi_req_wen0_i),
    .waddr1_i(mi_req_waddr1_i[8:0]),
    .wdata1_i(mi_req_wdata1_i[143:0]),
    .wen1_i(mi_req_wen1_i),
    .raddr0_i(mi_req_raddr0_i[8:0]),
    .rdata0_o(mi_req_rdata0_o[143:0]),
    .ren0_i(mi_req_ren0_i),
    .raddr1_i(mi_req_raddr1_i[8:0]),
    .rdata1_o(mi_req_rdata1_o[143:0]),
    .ren1_i(mi_req_ren1_i),
    .err_cor_o(mi_req_err_cor_o[5:0]),
    .err_uncor_o(mi_req_err_uncor_o[5:0])

  );

  generate 

  if (TL_COMPLETION_RAM_SIZE == 2'b10) begin : RAM32K

    xp4_usp_smsw_bram_32k #(

      .TCQ (TCQ),
      .TO_RAM_WRITE_PIPELINE(TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE),
      .TO_RAM_READ_PIPELINE(TL_RX_COMPLETION_TO_RAM_READ_PIPELINE),
      .FROM_RAM_READ_PIPELINE(TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE)

    )
    bram_comp_inst (

      .clk_i (core_clk_i),
      .reset_i (reset_i),
  
      .waddr0_i(mi_cpl_waddr0_i[8:0]),
      .wdata0_i(mi_cpl_wdata0_i[143:0]),
      .wen0_i(mi_cpl_wen0_i[1:0]),
      .waddr1_i(mi_cpl_waddr1_i[8:0]),
      .wdata1_i(mi_cpl_wdata1_i[143:0]),
      .wen1_i(mi_cpl_wen1_i[1:0]),
      .raddr0_i(mi_cpl_raddr0_i[8:0]),
      .rdata0_o(mi_cpl_rdata0_o[143:0]),
      .ren0_i(mi_cpl_ren0_i[1:0]),
      .raddr1_i(mi_cpl_raddr1_i[8:0]),
      .rdata1_o(mi_cpl_rdata1_o[143:0]),
      .ren1_i(mi_cpl_ren1_i[1:0]),
      .err_cor_o(mi_cpl_err_cor_o[11:0]),
      .err_uncor_o(mi_cpl_err_uncor_o[11:0])

    );

  end else begin : RAM16K

    xp4_usp_smsw_bram_16k #(

      .TCQ (TCQ),
      .TO_RAM_WRITE_PIPELINE(TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE),
      .TO_RAM_READ_PIPELINE(TL_RX_COMPLETION_TO_RAM_READ_PIPELINE),
      .FROM_RAM_READ_PIPELINE(TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE)

    )
    bram_comp_inst (

      .clk_i (core_clk_i),
      .reset_i (reset_i),
  
      .waddr0_i(mi_cpl_waddr0_i[8:0]),
      .wdata0_i(mi_cpl_wdata0_i[143:0]),
      .wen0_i(mi_cpl_wen0_i[0]),
      .waddr1_i(mi_cpl_waddr1_i[8:0]),
      .wdata1_i(mi_cpl_wdata1_i[143:0]),
      .wen1_i(mi_cpl_wen1_i[0]),
      .raddr0_i(mi_cpl_raddr0_i[8:0]),
      .rdata0_o(mi_cpl_rdata0_o[143:0]),
      .ren0_i(mi_cpl_ren0_i[0]),
      .raddr1_i(mi_cpl_raddr1_i[8:0]),
      .rdata1_o(mi_cpl_rdata1_o[143:0]),
      .ren1_i(mi_cpl_ren1_i[0]),
      .err_cor_o(mi_cpl_err_cor_o[5:0]),
      .err_uncor_o(mi_cpl_err_uncor_o[5:0])

    );

    assign mi_cpl_err_cor_o[11:6] = 6'b0;
    assign mi_cpl_err_uncor_o[11:6] = 6'b0;

  end

  endgenerate 

  xp4_usp_smsw_bram_msix #(

    .TCQ (TCQ),
    .TO_RAM_PIPELINE(AXISTEN_IF_MSIX_TO_RAM_PIPELINE),
    .FROM_RAM_PIPELINE(AXISTEN_IF_MSIX_FROM_RAM_PIPELINE),
    .MSIX_CAP_TABLE_SIZE(MSIX_CAP_TABLE_SIZE),
    .MSIX_TABLE_RAM_ENABLE(MSIX_TABLE_RAM_ENABLE)

  )
  bram_msix_inst (

    .clk_i(user_clk_i),
    .reset_i(reset_i),

    .addr_i(cfg_msix_waddr_i[12:0]),
    .wdata_i(cfg_msix_wdata_i[31:0]),
    .wdip_i(cfg_msix_wdip_i[3:0]),
    .wen_i(cfg_msix_wen_i[3:0]),
    .rdata_o(cfg_msix_rdata_o[31:0]),
    .rdop_o(cfg_msix_rdop_o[3:0])

  );

  xp4_usp_smsw_bram_tph #(

    .TCQ (TCQ),
    .TO_RAM_PIPELINE(TPH_TO_RAM_PIPELINE),
    .FROM_RAM_PIPELINE(TPH_FROM_RAM_PIPELINE),
    .TL_PF_ENABLE_REG(TL_PF_ENABLE_REG),
    .SRIOV_CAP_ENABLE(SRIOV_CAP_ENABLE),
    .PF0_SRIOV_CAP_TOTAL_VF(PF0_SRIOV_CAP_TOTAL_VF),
    .PF1_SRIOV_CAP_TOTAL_VF(PF1_SRIOV_CAP_TOTAL_VF),
    .PF2_SRIOV_CAP_TOTAL_VF(PF2_SRIOV_CAP_TOTAL_VF),
    .PF3_SRIOV_CAP_TOTAL_VF(PF3_SRIOV_CAP_TOTAL_VF),
    .PF0_TPHR_CAP_ENABLE(PF0_TPHR_CAP_ENABLE)

  )
  bram_tph_inst (

    .clk_i(user_clk_i),
    .reset_i(reset_i),

    .user_tph_stt_func_num_i(user_tph_stt_func_num_i[7:0]),
    .user_tph_stt_index_i(user_tph_stt_index_i[5:0]),
    .user_tph_stt_rd_en_i(user_tph_stt_rd_en_i),
    .user_tph_stt_rd_data_o(user_tph_stt_rd_data_o[7:0]),

    .addr_i(cfg_tph_waddr_i[11:0]),
    .wdata_i(cfg_tph_wdata_i[31:0]),
    .wdip_i(cfg_tph_wdip_i[3:0]),
    .wen_i(cfg_tph_wen_i[3:0]),
    .rdata_o(cfg_tph_rdata_o[31:0]),
    .rdop_o(cfg_tph_rdop_o[3:0])

  );

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_bram_16k_int.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_bram_16k_int #(

  parameter TCQ = 100

  ) (

  input  wire         clk_i,
  input  wire         reset_i,

  input  wire   [8:0] waddr0_i,
  input  wire   [0:0] wen0_i,
  input  wire [143:0] wdata0_i,
  input  wire   [8:0] waddr1_i,
  input  wire   [0:0] wen1_i,
  input  wire [143:0] wdata1_i,

  input  wire   [8:0] raddr0_i,
  input  wire   [0:0] ren0_i,
  output wire [143:0] rdata0_o,
  input  wire   [8:0] raddr1_i,
  input  wire   [0:0] ren1_i,
  output wire [143:0] rdata1_o,

  output wire   [5:0] err_cor_o,
  output wire   [5:0] err_uncor_o

  );

  genvar              i;

  wire [383:0]        rdata_w;
  wire [383:0]        wdata_w = {48'b0, wdata1_i[143:0], 48'b0, wdata0_i};

  generate begin : ECC_RAM

   for (i = 0; i < 6; i = i + 1)
   begin : RAMB36E2
        RAMB36E2 #(
          .DOA_REG (1),
          .DOB_REG (1),
          .EN_ECC_READ ("TRUE"),
          .EN_ECC_WRITE ("TRUE"),
          .INIT_A (36'h000000000),
          .INIT_B (36'h000000000),
          .INIT_FILE ("NONE"),
          .READ_WIDTH_A (72),
          .READ_WIDTH_B (0),
          .RSTREG_PRIORITY_A ("REGCE"),
          .RSTREG_PRIORITY_B ("REGCE"),
          .SIM_COLLISION_CHECK("ALL"),
          .SRVAL_A (36'h000000000),
          .SRVAL_B (36'h000000000),
          .WRITE_MODE_A ("WRITE_FIRST"),
          .WRITE_MODE_B ("WRITE_FIRST"),
          .WRITE_WIDTH_A (0),
          .WRITE_WIDTH_B (72))
        ramb36e2_inst (
          .ADDRENA (1'b1),
          .ADDRENB (1'b1),
          .CASDIMUXA (1'b0),
          .CASDIMUXB (1'b0),
          .CASDOMUXA (1'b0),
          .CASDOMUXB (1'b0),
          .CASDOMUXEN_A (1'b0),
          .CASDOMUXEN_B (1'b0),
          .CASINDBITERR (1'b0),
          .CASINSBITERR (1'b0),
          .CASOREGIMUXA (1'b0),
          .CASOREGIMUXB (1'b0),
          .CASOREGIMUXEN_A (1'b0),
          .CASOREGIMUXEN_B (1'b0),
          .ECCPIPECE (1'b0),
          .SLEEP (1'b0),
          .CASDINA (32'b0),
          .CASDINB (32'b0),
          .CASDINPA(4'b0),
          .CASDINPB(4'b0),
          .CASDOUTA (),
          .CASDOUTB (),
          .CASDOUTPA (),
          .CASDOUTPB (),
          .CASOUTDBITERR (),
          .CASOUTSBITERR (),
          .CLKARDCLK (clk_i),
          .CLKBWRCLK (clk_i),
          .DBITERR (err_uncor_o[i]),
          .ENARDEN ((i > 2) ? ren1_i : ren0_i),
          .ENBWREN ((i > 2) ? wen1_i : wen0_i),
          .INJECTDBITERR (1'b0),
          .INJECTSBITERR (1'b0),
          .REGCEAREGCE (1'b1),
          .REGCEB (1'b0),
          .RSTRAMARSTRAM (1'b0),
          .RSTRAMB (1'b0),
          .RSTREGARSTREG (1'b0),
          .RSTREGB (1'b0),
          .SBITERR (err_cor_o[i]),
          .ADDRARDADDR ({(i>2) ? raddr1_i[8:0] : raddr0_i[8:0], 6'b0}),
          .ADDRBWRADDR ({(i>2) ? waddr1_i[8:0] : waddr0_i[8:0], 6'b0}),
          .DINADIN (wdata_w[(2*32*i)+31:(2*32*i)+0]),
          .DINBDIN (wdata_w[(2*32*i)+63:(2*32*i)+32]),
          .DINPADINP (4'b0),
          .DINPBDINP (4'b0),
          .DOUTADOUT (rdata_w[(2*32*i)+31:(2*32*i)+0]),
          .DOUTBDOUT (rdata_w[(2*32*i)+63:(2*32*i)+32]),
          .DOUTPADOUTP (),
          .DOUTPBDOUTP (),
          .ECCPARITY (),
          .RDADDRECC (),
          .WEA (4'h0),
          .WEBWE (8'hFF)
        );
      end
    end
  endgenerate

  assign rdata1_o =  rdata_w[335:192];
  assign rdata0_o =  rdata_w[143:000];

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_bram_16k.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_bram_16k #(

  parameter           TCQ = 100
, parameter           TO_RAM_WRITE_PIPELINE="FALSE"
, parameter           TO_RAM_READ_PIPELINE="FALSE"
, parameter           FROM_RAM_READ_PIPELINE="FALSE"

  ) (

  input  wire         clk_i,
  input  wire         reset_i,

  input  wire   [8:0] waddr0_i,
  input  wire   [0:0] wen0_i,
  input  wire [143:0] wdata0_i,
  input  wire   [8:0] waddr1_i,
  input  wire   [0:0] wen1_i,
  input  wire [143:0] wdata1_i,

  input  wire   [8:0] raddr0_i,
  input  wire   [0:0] ren0_i,
  output wire [143:0] rdata0_o,
  input  wire   [8:0] raddr1_i,
  input  wire   [0:0] ren1_i,
  output wire [143:0] rdata1_o,

  output wire   [5:0] err_cor_o,
  output wire   [5:0] err_uncor_o

  );

  reg           [8:0] waddr0;
  reg           [0:0] wen0;
  reg         [143:0] wdata0;
  reg           [8:0] waddr1;
  reg           [0:0] wen1;
  reg         [143:0] wdata1;
  reg           [8:0] raddr0;
  reg           [0:0] ren0;
  reg           [8:0] raddr1;
  reg           [0:0] ren1;
  wire        [143:0] rdata0;
  wire        [143:0] rdata1;
  wire          [5:0] err_cor;
  wire          [5:0] err_uncor;
  reg         [143:0] reg_rdata0;
  reg         [143:0] reg_rdata1;
  reg           [5:0] reg_err_cor;
  reg           [5:0] reg_err_uncor;

  //
  // Optional input pipe stages
  //
  generate

    if (TO_RAM_WRITE_PIPELINE == "TRUE") begin : TOWRPIPELINE

      always @(posedge clk_i) begin
     
        if (reset_i) begin

          waddr0 <= #(TCQ) 9'b0;
          wen0 <= #(TCQ) 1'b0;
          wdata0 <= #(TCQ) 144'b0;
          waddr1 <= #(TCQ) 9'b0;
          wen1 <= #(TCQ) 1'b0;
          wdata1 <= #(TCQ) 144'b0;

        end else begin

          waddr0 <= #(TCQ) waddr0_i;
          wen0 <= #(TCQ) wen0_i;
          wdata0 <= #(TCQ) wdata0_i;
          waddr1 <= #(TCQ) waddr1_i;
          wen1 <= #(TCQ) wen1_i;
          wdata1 <= #(TCQ) wdata1_i;

        end

      end

    end else begin : NOTOWRPIPELINE

      always @(*) begin

        waddr0 = waddr0_i;
        wen0 = wen0_i;
        wdata0 = wdata0_i;
        waddr1 = waddr1_i;
        wen1 = wen1_i;
        wdata1 = wdata1_i;

      end

    end

    if (TO_RAM_READ_PIPELINE == "TRUE") begin : TORDPIPELINE

      always @(posedge clk_i) begin
     
        if (reset_i) begin

          raddr0 <= #(TCQ) 9'b0;
          ren0 <= #(TCQ) 1'b0;
          raddr1 <= #(TCQ) 9'b0;
          ren1 <= #(TCQ) 1'b0;

        end else begin

          raddr0 <= #(TCQ) raddr0_i;
          ren0 <= #(TCQ) ren0_i;
          raddr1 <= #(TCQ) raddr1_i;
          ren1 <= #(TCQ) ren1_i;

        end

      end

    end else begin : NOTORDPIPELINE

      always @(*) begin

        raddr0 = raddr0_i;
        ren0 = ren0_i;
        raddr1 = raddr1_i;
        ren1 = ren1_i;

      end

    end
  
  endgenerate

  //
  // Optional output pipe stages
  //
  generate

    if (FROM_RAM_READ_PIPELINE == "TRUE") begin : FRMRDPIPELINE


      always @(posedge clk_i) begin
     
        if (reset_i) begin

          reg_rdata0 <= #(TCQ) 144'b0;
          reg_rdata1 <= #(TCQ) 144'b0;
          reg_err_cor <= #(TCQ) 6'b0;
          reg_err_uncor <= #(TCQ) 6'b0;

         end else begin

          reg_rdata0 <= #(TCQ) rdata0;
          reg_rdata1 <= #(TCQ) rdata1;
          reg_err_cor <= #(TCQ) err_cor;
          reg_err_uncor <= #(TCQ) err_uncor;

        end

      end

    end else begin : NOFRMRDPIPELINE

      always @(*) begin

          reg_rdata0 = rdata0;
          reg_rdata1 = rdata1;
          reg_err_cor = err_cor;
          reg_err_uncor = err_uncor;

      end

    end
  
  endgenerate

  assign rdata0_o = reg_rdata0;
  assign rdata1_o = reg_rdata1;
  assign err_cor_o = reg_err_cor;
  assign err_uncor_o = reg_err_uncor;

  xp4_usp_smsw_bram_16k_int #(
      .TCQ(TCQ)
    )
    bram_16k_int (

      .clk_i (clk_i),
      .reset_i (reset_i),

      .waddr0_i(waddr0[8:0]),
      .wdata0_i(wdata0[143:0]),
      .wen0_i(wen0),
      .waddr1_i(waddr1[8:0]),
      .wdata1_i(wdata1[143:0]),
      .wen1_i(wen1),
      .raddr0_i(raddr0[8:0]),
      .rdata0_o(rdata0[143:0]),
      .ren0_i(ren0),
      .raddr1_i(raddr1[8:0]),
      .rdata1_o(rdata1[143:0]),
      .ren1_i(ren1),
      .err_cor_o(err_cor[5:0]),
      .err_uncor_o(err_uncor[5:0])

  );


endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_bram_32k.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_bram_32k #(

  parameter           TCQ = 100
, parameter           TO_RAM_WRITE_PIPELINE="FALSE"
, parameter           TO_RAM_READ_PIPELINE="FALSE"
, parameter           FROM_RAM_READ_PIPELINE="FALSE"

  ) (

  input  wire         clk_i,
  input  wire         reset_i,

  input  wire   [8:0] waddr0_i,
  input  wire   [1:0] wen0_i,
  input  wire [143:0] wdata0_i,
  input  wire   [8:0] waddr1_i,
  input  wire   [1:0] wen1_i,
  input  wire [143:0] wdata1_i,

  input  wire   [8:0] raddr0_i,
  input  wire   [1:0] ren0_i,
  output wire [143:0] rdata0_o,
  input  wire   [8:0] raddr1_i,
  input  wire   [1:0] ren1_i,
  output wire [143:0] rdata1_o,

  output wire   [11:0] err_cor_o,
  output wire   [11:0] err_uncor_o

  );

  wire [143:0] rdata0_0;
  wire [143:0] rdata0_1;
  wire [143:0] rdata1_0;
  wire [143:0] rdata1_1;

  wire  [11:0] err_cor;
  wire  [11:0] err_uncor;

  reg  [143:0] reg_rdata0;
  reg  [143:0] reg_rdata1;
  reg   [11:0] reg_err_cor;
  reg   [11:0] reg_err_uncor;

  reg    [0:0] reg_raddr0_10_p0;
  reg    [0:0] reg_raddr1_10_p0;
  (* keep = "true", max_fanout = 32 *) reg    [0:0] reg_raddr0_10_p1;
  (* keep = "true", max_fanout = 32 *) reg    [0:0] reg_raddr1_10_p1;
  wire   [0:0] raddr0_10_p0;
  wire   [0:0] raddr1_10_p0;

  reg    [8:0] raddr0;
  reg    [1:0] ren0;
  reg    [8:0] raddr1;
  reg    [1:0] ren1;

  reg    [8:0] waddr0;
  reg    [1:0] wen0;
  reg  [143:0] wdata0;
  reg    [8:0] waddr1;
  reg    [1:0] wen1;
  reg  [143:0] wdata1;
  
  //
  // Optional input pipe stages
  //
  generate

    if (TO_RAM_WRITE_PIPELINE == "TRUE") begin : TOWRPIPELINE

      always @(posedge clk_i) begin
     
        if (reset_i) begin

          waddr0 <= #(TCQ) 9'b0;
          wen0 <= #(TCQ) 2'b0;
          wdata0 <= #(TCQ) 144'b0;
          waddr1 <= #(TCQ) 9'b0;
          wen1 <= #(TCQ) 2'b0;
          wdata1 <= #(TCQ) 144'b0;

	end else begin

          waddr0 <= #(TCQ) waddr0_i;
          wen0 <= #(TCQ) wen0_i;
          wdata0 <= #(TCQ) wdata0_i;
          waddr1 <= #(TCQ) waddr1_i;
          wen1 <= #(TCQ) wen1_i;
          wdata1 <= #(TCQ) wdata1_i;

	end

     end

    end else begin : NOTOWRPIPELINE

      always @(*) begin

        waddr0 = waddr0_i;
        wen0 = wen0_i;
        wdata0 = wdata0_i;
        waddr1 = waddr1_i;
        wen1 = wen1_i;
        wdata1 = wdata1_i;
    
      end
  
    end

    if (TO_RAM_READ_PIPELINE == "TRUE") begin : TORDPIPELINE

      always @(posedge clk_i) begin
     
        if (reset_i) begin

          raddr0 <= #(TCQ) 9'b0;
          ren0 <= #(TCQ) 1'b0;
          raddr1 <= #(TCQ) 9'b0;
          ren1 <= #(TCQ) 1'b0;

	end else begin

          raddr0 <= #(TCQ) raddr0_i;
          ren0 <= #(TCQ) ren0_i;
          raddr1 <= #(TCQ) raddr1_i;
          ren1 <= #(TCQ) ren1_i;

	end

      end

    end else begin : NOTORDPIPELINE

      always @(*) begin

        raddr0 = raddr0_i;
        ren0 = ren0_i;
        raddr1 = raddr1_i;
        ren1 = ren1_i;

      end

    end
  
  endgenerate
 
  //
  // output pipe stage
  //

  generate

    if (FROM_RAM_READ_PIPELINE == "TRUE") begin : FRMRDPIPELINE

      always @(posedge clk_i) begin
     
        if (reset_i) begin

          reg_rdata0 <= #(TCQ) 144'b0;
          reg_rdata1 <= #(TCQ) 144'b0;
          reg_err_cor <= #(TCQ) 12'b0;
          reg_err_uncor <= #(TCQ) 12'b0;
    
        end else begin
    
          reg_rdata0 <= #(TCQ) raddr0_10_p0 ? rdata1_0 : rdata0_0;
          reg_rdata1 <= #(TCQ) raddr1_10_p0 ? rdata1_1 : rdata0_1;
          reg_err_cor <= #(TCQ) err_cor;
          reg_err_uncor <= #(TCQ) err_uncor;
    
        end
    
      end

   end else begin : NOFRMRDPIPELINE

      always @(*) begin

        reg_rdata0 = raddr0_10_p0 ? rdata1_0 : rdata0_0;
        reg_rdata1 = raddr1_10_p0 ? rdata1_1 : rdata0_1;
        reg_err_cor = err_cor;
        reg_err_uncor = err_uncor;

      end

   end

  endgenerate

  always @(posedge clk_i) begin
     
    if (reset_i) begin

      reg_raddr0_10_p0 <= #(TCQ) 1'b0;
      reg_raddr1_10_p0 <= #(TCQ) 1'b0;
      reg_raddr0_10_p1 <= #(TCQ) 1'b0;
      reg_raddr1_10_p1 <= #(TCQ) 1'b0;
    
    end else begin
    
      reg_raddr0_10_p0 <= #(TCQ) ren0[1];
      reg_raddr1_10_p0 <= #(TCQ) ren1[1];
      reg_raddr0_10_p1 <= #(TCQ) reg_raddr0_10_p0;
      reg_raddr1_10_p1 <= #(TCQ) reg_raddr1_10_p0;
    
    end
    
  end

  assign rdata0_o = reg_rdata0;
  assign rdata1_o = reg_rdata1;
  assign err_cor_o = reg_err_cor;
  assign err_uncor_o = reg_err_uncor;
  assign raddr0_10_p0 = reg_raddr0_10_p1;
  assign raddr1_10_p0 = reg_raddr1_10_p1;

  // Upper 512 Words
  xp4_usp_smsw_bram_16k_int #( 
	.TCQ(TCQ)) 
  bram_16k_0_int (
    .clk_i (clk_i),
    .reset_i (reset_i),

    .waddr0_i(waddr0[8:0]),
    .wdata0_i(wdata0[143:0]),
    .wen0_i(wen0[0]),
    .waddr1_i(waddr1[8:0]),
    .wdata1_i(wdata1[143:0]),
    .wen1_i(wen1[0]),
    .raddr0_i(raddr0[8:0]),
    .rdata0_o(rdata0_0[143:0]),
    .ren0_i(ren0[0]),
    .raddr1_i(raddr1[8:0]),
    .rdata1_o(rdata0_1[143:0]),
    .ren1_i(ren1[0]),
    .err_cor_o(err_cor[5:0]),
    .err_uncor_o(err_uncor[5:0])

  );
  
  // Lower 512 Words
  xp4_usp_smsw_bram_16k_int #( 
	.TCQ(TCQ)) 
  bram_16k_1_int (
    .clk_i (clk_i),
    .reset_i (reset_i),

    .waddr0_i(waddr0[8:0]),
    .wdata0_i(wdata0[143:0]),
    .wen0_i(wen0[1]),
    .waddr1_i(waddr1[8:0]),
    .wdata1_i(wdata1[143:0]),
    .wen1_i(wen1[1]),
    .raddr0_i(raddr0[8:0]),
    .rdata0_o(rdata1_0[143:0]),
    .ren0_i(ren0[1]),
    .raddr1_i(raddr1[8:0]),
    .rdata1_o(rdata1_1[143:0]),
    .ren1_i(ren1[1]),
    .err_cor_o(err_cor[11:6]),
    .err_uncor_o(err_uncor[11:6])

  );

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_bram_4k_int.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_bram_4k_int #(
  parameter TCQ = 100
  ) (
  input  wire         clk_i,
  input  wire         reset_i,
  input  wire   [9:0] addr_i,
  input  wire  [31:0] wdata_i,
  input  wire   [3:0] wdip_i,
  input  wire   [3:0] wen_i,
  output wire  [31:0] rdata_o,
  output wire   [3:0] rdop_o,
  input  wire   [9:0] baddr_i,
  output wire  [31:0] brdata_o
  );

  genvar              i;

  RAMB36E2 #(
        .DOA_REG (1),
        .DOB_REG (1),
        .EN_ECC_READ ("FALSE"),
        .EN_ECC_WRITE ("FALSE"),
        .INIT_A (36'h000000000),
        .INIT_B (36'h000000000),
        .INIT_FILE ("NONE"),
        .READ_WIDTH_A (36),
        .READ_WIDTH_B (36),
        .RSTREG_PRIORITY_A ("REGCE"),
        .RSTREG_PRIORITY_B ("REGCE"),
        .SIM_COLLISION_CHECK("GENERATE_X_ONLY"),
        .SRVAL_A (36'h000000000),
        .SRVAL_B (36'h000000000),
        .WRITE_MODE_A ("WRITE_FIRST"),
        .WRITE_MODE_B ("WRITE_FIRST"),
        .WRITE_WIDTH_A (36),
        .WRITE_WIDTH_B (36))
  ramb36e2_inst (
        .ADDRENA (1'b1),
        .ADDRENB (1'b1),
        .CASDIMUXA (1'b0),
        .CASDIMUXB (1'b0),
        .CASDOMUXA (1'b0),
        .CASDOMUXB (1'b0),
        .CASDOMUXEN_A (1'b0),
        .CASDOMUXEN_B (1'b0),
        .CASINDBITERR (1'b0),
        .CASINSBITERR (1'b0),
        .CASOREGIMUXA (1'b0),
        .CASOREGIMUXB (1'b0),
        .CASOREGIMUXEN_A (1'b0),
        .CASOREGIMUXEN_B (1'b0),
        .ECCPIPECE (1'b0),
        .SLEEP (1'b0),
        .CASDINA (32'b0),
        .CASDINB (32'b0),
        .CASDINPA(4'b0),
        .CASDINPB(4'b0),
        .CASDOUTA (),
        .CASDOUTB (),
        .CASDOUTPA (),
        .CASDOUTPB (),
        .CASOUTDBITERR (),
        .CASOUTSBITERR (),
        .CLKARDCLK (clk_i),
        .CLKBWRCLK (clk_i),
        .DBITERR (),
        .ENARDEN (1'b1),
        .ENBWREN (1'b1),
        .INJECTDBITERR (1'b0),
        .INJECTSBITERR (1'b0),
        .REGCEAREGCE (1'b1),
        .REGCEB (1'b1),
        .RSTRAMARSTRAM (1'b0),
        .RSTRAMB (1'b0),
        .RSTREGARSTREG (1'b0),
        .RSTREGB (1'b0),
        .SBITERR (),
        .ADDRARDADDR ({addr_i[9:0], 5'b0}),
        .ADDRBWRADDR ({baddr_i[9:0], 5'b0}),
        .DINADIN (wdata_i[31:0]),
        .DINBDIN (32'b0),
        .DINPADINP (wdip_i[3:0]),
        .DINPBDINP (4'b0),
        .DOUTADOUT (rdata_o[31:0]),
        .DOUTBDOUT (brdata_o[31:0]),
        .DOUTPADOUTP (rdop_o[3:0]),
        .DOUTPBDOUTP (),
        .ECCPARITY (),
        .RDADDRECC (),
        .WEA (wen_i[3:0]),
        .WEBWE (8'b0)
      );

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_bram_msix.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_bram_msix #(

  parameter           TCQ = 100
, parameter           TO_RAM_PIPELINE="FALSE"
, parameter           FROM_RAM_PIPELINE="FALSE"
, parameter           MSIX_CAP_TABLE_SIZE=11'h0
, parameter           MSIX_TABLE_RAM_ENABLE="FALSE"

  ) (

  input  wire         clk_i,
  input  wire         reset_i,

  input  wire  [12:0] addr_i,
  input  wire  [31:0] wdata_i,
  input  wire   [3:0] wdip_i,
  input  wire   [3:0] wen_i,
  output wire  [31:0] rdata_o,
  output wire   [3:0] rdop_o

  );

  // WIP : Use Total number of functions (PFs + VFs) to calculate the NUM_BRAM_4K
  localparam integer NUM_BRAM_4K = (MSIX_TABLE_RAM_ENABLE == "TRUE") ? 8 : 0 ;
 

  reg          [12:0] addr;
  reg          [12:0] addr_p0;
  reg          [12:0] addr_p1;
  reg          [31:0] wdata;
  reg           [3:0] wdip;
  reg           [3:0] wen;
  reg          [31:0] reg_rdata;
  reg           [3:0] reg_rdop;
  wire         [31:0] rdata;
  wire          [3:0] rdop;
  genvar              i;
  wire    [(8*4)-1:0] bram_4k_wen;
  wire   [(8*32)-1:0] rdata_t;
  wire    [(8*4)-1:0] rdop_t;

  //
  // Optional input pipe stages
  //
  generate

    if (TO_RAM_PIPELINE == "TRUE") begin : TORAMPIPELINE

      always @(posedge clk_i) begin
     
        if (reset_i) begin

          addr <= #(TCQ) 13'b0;
          wdata <= #(TCQ) 32'b0;
          wdip <= #(TCQ) 4'b0;
          wen <= #(TCQ) 4'b0;

        end else begin

          addr <= #(TCQ) addr_i;
          wdata <= #(TCQ) wdata_i;
          wdip <= #(TCQ) wdip_i;
          wen <= #(TCQ) wen_i;

        end

      end

    end else begin : NOTORAMPIPELINE

      always @(*) begin

          addr = addr_i;
          wdata = wdata_i;
          wdip = wdip_i;
          wen = wen_i;

      end


    end

  endgenerate

  // 
  // Address pipeline
  //
  always @(posedge clk_i) begin
     
    if (reset_i) begin

      addr_p0 <= #(TCQ) 13'b0;
      addr_p1 <= #(TCQ) 13'b0;

    end else begin

      addr_p0 <= #(TCQ) addr;
      addr_p1 <= #(TCQ) addr_p0;

    end

  end

  //
  // Optional output pipe stages
  //
  generate

    if (FROM_RAM_PIPELINE == "TRUE") begin : FRMRAMPIPELINE


      always @(posedge clk_i) begin
     
        if (reset_i) begin

          reg_rdata <= #(TCQ) 32'b0;
          reg_rdop <= #(TCQ) 4'b0;

        end else begin

          case (addr_p1[12:10]) 
            3'b000 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(0))+31:(32*(0))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(0))+3:(4*(0))+0];
            end
            3'b001 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(1))+31:(32*(1))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(1))+3:(4*(1))+0];
            end
            3'b010 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(2))+31:(32*(2))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(2))+3:(4*(2))+0];
            end
            3'b011 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(3))+31:(32*(3))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(3))+3:(4*(3))+0];
            end
            3'b100 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(4))+31:(32*(4))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(4))+3:(4*(4))+0];
            end
            3'b101 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(5))+31:(32*(5))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(5))+3:(4*(5))+0];
            end
            3'b110 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(6))+31:(32*(6))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(6))+3:(4*(6))+0];
            end
            3'b111 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(7))+31:(32*(7))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(7))+3:(4*(7))+0];
            end
          endcase

        end

      end

    end else begin : NOFRMRAMPIPELINE

      always @(*) begin

          case (addr_p1[12:10]) 
            3'b000 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(0))+31:(32*(0))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(0))+3:(4*(0))+0];
            end
            3'b001 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(1))+31:(32*(1))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(1))+3:(4*(1))+0];
            end
            3'b010 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(2))+31:(32*(2))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(2))+3:(4*(2))+0];
            end
            3'b011 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(3))+31:(32*(3))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(3))+3:(4*(3))+0];
            end
            3'b100 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(4))+31:(32*(4))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(4))+3:(4*(4))+0];
            end
            3'b101 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(5))+31:(32*(5))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(5))+3:(4*(5))+0];
            end
            3'b110 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(6))+31:(32*(6))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(6))+3:(4*(6))+0];
            end
            3'b111 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(7))+31:(32*(7))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(7))+3:(4*(7))+0];
            end
          endcase

      end

    end
  
  endgenerate

  assign rdata_o = (MSIX_TABLE_RAM_ENABLE == "TRUE") ?  reg_rdata : 32'h0;
  assign rdop_o = (MSIX_TABLE_RAM_ENABLE == "TRUE") ? reg_rdop : 4'h0;

  generate 
  
    for (i=0; i<NUM_BRAM_4K; i=i+1) begin : BRAM4K

      xp4_usp_smsw_bram_4k_int #(
          .TCQ(TCQ)
        )
        bram_4k_int (
    
          .clk_i (clk_i),
          .reset_i (reset_i),
    
          .addr_i(addr[9:0]),
          .wdata_i(wdata),
          .wdip_i(wdip),
          .wen_i(bram_4k_wen[(4*(i))+3:(4*(i))+0]),
          .rdata_o(rdata_t[(32*i)+31:(32*i)+0]),
          .rdop_o(rdop_t[(4*i)+3:(4*i)+0]),
          .baddr_i(10'b0),
          .brdata_o()

      );
      assign bram_4k_wen[(4*(i))+3:(4*(i))+0] = wen & {4{(i == addr[12:10])}};  
      
    end

  endgenerate

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_bram_rep_int.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_bram_rep_int #(

  parameter TCQ = 100

  ) (

  input  wire         clk_i,
  input  wire         reset_i,

  input  wire   [8:0] addr_i,
  input  wire   [0:0] wen_i,
  input  wire [255:0] wdata_i,
  input  wire   [0:0] ren_i,
  output wire [255:0] rdata_o,

  output wire   [3:0] err_cor_o,
  output wire   [3:0] err_uncor_o

  );

  genvar              i;

  wire [255:0]        rdata_w;
  wire [255:0]        wdata_w = wdata_i;

  generate begin : ECC_RAM

   for (i = 0; i < 4; i = i + 1)
   begin : RAMB36E2
        RAMB36E2 #(
          .DOA_REG (1),
          .DOB_REG (1),
          .EN_ECC_READ ("TRUE"),
          .EN_ECC_WRITE ("TRUE"),
          .INIT_A (36'h000000000),
          .INIT_B (36'h000000000),
          .INIT_FILE ("NONE"),
          .READ_WIDTH_A (72),
          .READ_WIDTH_B (0),
          .RSTREG_PRIORITY_A ("REGCE"),
          .RSTREG_PRIORITY_B ("REGCE"),
          .SIM_COLLISION_CHECK ("ALL"),
          .SRVAL_A (36'h000000000),
          .SRVAL_B (36'h000000000),
          .WRITE_MODE_A ("WRITE_FIRST"),
          .WRITE_MODE_B ("WRITE_FIRST"),
          .WRITE_WIDTH_A (0),
          .WRITE_WIDTH_B (72))
        ramb36e2_inst (
          .ADDRENA (1'b1),
          .ADDRENB (1'b1),
          .CASDIMUXA (1'b0),
          .CASDIMUXB (1'b0),
          .CASDOMUXA (1'b0),
          .CASDOMUXB (1'b0),
          .CASDOMUXEN_A (1'b0),
          .CASDOMUXEN_B (1'b0),
          .CASINDBITERR (1'b0),
          .CASINSBITERR (1'b0),
          .CASOREGIMUXA (1'b0),
          .CASOREGIMUXB (1'b0),
          .CASOREGIMUXEN_A (1'b0),
          .CASOREGIMUXEN_B (1'b0),
          .ECCPIPECE (1'b0),
          .SLEEP (1'b0),
          .CASDINA (32'b0),
          .CASDINB (32'b0),
          .CASDINPA(4'b0),
          .CASDINPB(4'b0),
          .CASDOUTA (),
          .CASDOUTB (),
          .CASDOUTPA (),
          .CASDOUTPB (),
          .CASOUTDBITERR (),
          .CASOUTSBITERR (),
          .CLKARDCLK (clk_i),
          .CLKBWRCLK (clk_i),
          .DBITERR (err_uncor_o[i]),
          .ENARDEN (ren_i),
          .ENBWREN (wen_i),
          .INJECTDBITERR (1'b0),
          .INJECTSBITERR (1'b0),
          .REGCEAREGCE (1'b1),
          .REGCEB (1'b0),
          .RSTRAMARSTRAM (1'b0),
          .RSTRAMB (1'b0),
          .RSTREGARSTREG (1'b0),
          .RSTREGB (1'b0),
          .SBITERR (err_cor_o[i]),
          .ADDRARDADDR ({addr_i[8:0], 6'b0}),
          .ADDRBWRADDR ({addr_i[8:0], 6'b0}),
          .DINADIN (wdata_w[(2*32*i)+31:(2*32*i)+0]),
          .DINBDIN (wdata_w[(2*32*i)+63:(2*32*i)+32]),
          .DINPADINP (4'b0),
          .DINPBDINP (4'b0),
          .DOUTADOUT (rdata_w[(2*32*i)+31:(2*32*i)+0]),
          .DOUTBDOUT (rdata_w[(2*32*i)+63:(2*32*i)+32]),
          .DOUTPADOUTP (),
          .DOUTPBDOUTP (),
          .ECCPARITY (),
          .RDADDRECC (),
          .WEA (4'h0),
          .WEBWE (8'hFF)
        );
      end
    end
  endgenerate

  assign rdata_o =  rdata_w;

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_bram_rep.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_bram_rep #(
  parameter           TCQ = 100
, parameter           TO_RAM_PIPELINE="FALSE"
, parameter           FROM_RAM_PIPELINE="FALSE"

  ) (

  input  wire         clk_i,
  input  wire         reset_i,

  input  wire   [8:0] addr_i,
  input  wire   [0:0] wen_i,
  input  wire [255:0] wdata_i,

  output wire [255:0] rdata_o,
  input  wire   [0:0] ren_i,

  output wire   [3:0] err_cor_o,
  output wire   [3:0] err_uncor_o

  );

  reg           [8:0] addr;
  reg           [0:0] wen;
  reg           [0:0] ren;
  reg         [255:0] wdata;

  wire        [255:0] rdata;
  wire          [3:0] err_cor;
  wire          [3:0] err_uncor;

  reg         [255:0] reg_rdata;
  reg           [3:0] reg_err_cor;
  reg           [3:0] reg_err_uncor;

  //
  // Optional input pipe stages
  //
  
  generate

    if (TO_RAM_PIPELINE == "TRUE") begin : TORAMPIPELINE

      always @(posedge clk_i) begin
     
        if (reset_i) begin

          addr <= #(TCQ) 9'b0;
          wen <= #(TCQ) 1'b0;
          wdata <= #(TCQ) 256'b0;
          ren <= #(TCQ) 1'b0;

        end else begin

          addr <= #(TCQ) addr_i;
          wen <= #(TCQ) wen_i;
          wdata <= #(TCQ) wdata_i;
          ren <= #(TCQ) ren_i;

        end

      end

    end else begin : NOTORAMPIPELINE

      always @(*) begin

        addr = addr_i;
        wen = wen_i;
        wdata = wdata_i;
        ren = ren_i;

      end

    end

  endgenerate

  //
  // Optional output pipe stages
  //
  
  generate

    if (FROM_RAM_PIPELINE == "TRUE") begin : FRMRAMPIPELINE


      always @(posedge clk_i) begin
     
        if (reset_i) begin

          reg_rdata <= #(TCQ) 256'b0;
          reg_err_cor <= #(TCQ) 4'b0;
          reg_err_uncor <= #(TCQ) 4'b0;

        end else begin

          reg_rdata <= #(TCQ) rdata;
          reg_err_cor <= #(TCQ) err_cor;
          reg_err_uncor <= #(TCQ) err_uncor;

        end

      end

    end else begin : NOFRMRAMPIPELINE

      always @(*) begin

        reg_rdata = rdata;
        reg_err_cor = err_cor;
        reg_err_uncor = err_uncor;

      end

    end
  
  endgenerate

  assign rdata_o = reg_rdata;

  assign err_cor_o = reg_err_cor;
  assign err_uncor_o = reg_err_uncor;

  xp4_usp_smsw_bram_rep_int #(
      .TCQ(TCQ)
    )
    bram_rep_int_0 (

      .clk_i (clk_i),
      .reset_i (reset_i),

      .addr_i(addr[8:0]),
      .wdata_i(wdata[255:0]),
      .wen_i(wen),
      .ren_i(ren),
      .rdata_o(rdata[255:0]),
      .err_cor_o(err_cor[3:0]),
      .err_uncor_o(err_uncor[3:0])

  );


endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_bram_tph.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_bram_tph #(
  parameter           TCQ = 100
, parameter           TO_RAM_PIPELINE="FALSE"
, parameter           FROM_RAM_PIPELINE="FALSE"
, parameter [1:0]     TL_PF_ENABLE_REG=2'h0
, parameter [3:0]     SRIOV_CAP_ENABLE=4'h0
, parameter [15:0]    PF0_SRIOV_CAP_TOTAL_VF=16'h0
, parameter [15:0]    PF1_SRIOV_CAP_TOTAL_VF=16'h0
, parameter [15:0]    PF2_SRIOV_CAP_TOTAL_VF=16'h0
, parameter [15:0]    PF3_SRIOV_CAP_TOTAL_VF=16'h0
, parameter           PF0_TPHR_CAP_ENABLE="FALSE"

  ) (

  input  wire         clk_i,
  input  wire         reset_i,

  input  wire   [7:0] user_tph_stt_func_num_i,     // 0-255
  input  wire   [5:0] user_tph_stt_index_i,        // 0-63
  input  wire         user_tph_stt_rd_en_i,
  output wire   [7:0] user_tph_stt_rd_data_o,

  input  wire  [11:0] addr_i,
  input  wire  [31:0] wdata_i,
  input  wire   [3:0] wdip_i,
  input  wire   [3:0] wen_i,
  output wire  [31:0] rdata_o,
  output wire   [3:0] rdop_o

  );
  localparam integer NUM_VFUNCTIONS = (SRIOV_CAP_ENABLE == 4'h0) ? 0 : 
                              (SRIOV_CAP_ENABLE == 4'h1) ? PF0_SRIOV_CAP_TOTAL_VF : 
                              (SRIOV_CAP_ENABLE == 4'h3) ? (PF0_SRIOV_CAP_TOTAL_VF + PF1_SRIOV_CAP_TOTAL_VF) : 
                              (SRIOV_CAP_ENABLE == 4'h7) ? (PF0_SRIOV_CAP_TOTAL_VF + PF1_SRIOV_CAP_TOTAL_VF + PF2_SRIOV_CAP_TOTAL_VF) : 
                              (PF0_SRIOV_CAP_TOTAL_VF + PF1_SRIOV_CAP_TOTAL_VF + PF2_SRIOV_CAP_TOTAL_VF + PF3_SRIOV_CAP_TOTAL_VF);

  localparam integer NUM_FUNCTIONS = (TL_PF_ENABLE_REG == 2'h0) ? (NUM_VFUNCTIONS + 1) :
                             (TL_PF_ENABLE_REG == 2'h1) ? (NUM_VFUNCTIONS + 2) :
                             (TL_PF_ENABLE_REG == 2'h2) ? (NUM_VFUNCTIONS + 3) : (NUM_VFUNCTIONS + 4);

  localparam integer NUM_BRAM_4K = (PF0_TPHR_CAP_ENABLE == "TRUE") ?  
                                   ((NUM_FUNCTIONS  <= 64) ? 1 : 
                                   ((NUM_FUNCTIONS  > 64) && (NUM_FUNCTIONS  <= 128)) ? 2 : 
                                   ((NUM_FUNCTIONS  > 128) && (NUM_FUNCTIONS  <= 192)) ? 3 : 4) : 4;
 

  reg          [11:0] addr;
  reg          [11:0] addr_p0;
  reg          [11:0] addr_p1;
  reg          [31:0] wdata;
  reg           [3:0] wdip;
  reg           [3:0] wen;
  reg          [31:0] reg_rdata;
  reg           [3:0] reg_rdop;
  wire         [31:0] rdata;
  wire          [3:0] rdop;
  genvar              i;
  wire         [13:0] baddr; 
  reg          [13:0] baddr_p0; 
  reg          [13:0] baddr_p1; 
  reg          [31:0] brdata_w;
  wire   [(4*32)-1:0] rdata_t;
  wire    [(4*4)-1:0] rdop_t;
  wire   [(4*32)-1:0] brdata;
  wire    [(4*4)-1:0] bram_4k_wen;

  generate

    if (PF0_TPHR_CAP_ENABLE == "TRUE") begin : TPHR_CAP_PRESENT

      //
      // Optional input pipe stages
      //

      if (TO_RAM_PIPELINE == "TRUE") begin : TORAMPIPELINE

        always @(posedge clk_i) begin
     
          if (reset_i) begin

            addr <= #(TCQ) 12'b0;
            wdata <= #(TCQ) 32'b0;
            wdip <= #(TCQ) 4'b0;
            wen <= #(TCQ) 4'b0;
    
          end else begin
    
            addr <= #(TCQ) addr_i;
            wdata <= #(TCQ) wdata_i;
            wdip <= #(TCQ) wdip_i;
            wen <= #(TCQ) wen_i;
    
          end

        end

      end else begin : NOTORAMPIPELINE

        always @(*) begin

          addr = addr_i;
          wdata = wdata_i;
          wdip = wdip_i;
          wen = wen_i;
    
      end

    end


    // 
    // Address pipeline
    //

    always @(posedge clk_i) begin
     
      if (reset_i) begin

        addr_p0 <= #(TCQ) 12'b0;
        addr_p1 <= #(TCQ) 12'b0;
        baddr_p0 <= #(TCQ) 2'b0;
        baddr_p1 <= #(TCQ) 2'b0;
    
      end else begin
    
        addr_p0 <= #(TCQ) addr;
        addr_p1 <= #(TCQ) addr_p0;
        baddr_p0 <= #(TCQ) baddr;
        baddr_p1 <= #(TCQ) baddr_p0;
    
      end
    
    end

    //
    // Optional output pipe stages
    //

    if (FROM_RAM_PIPELINE == "TRUE") begin : FRMRAMPIPELINE
    
    
      always @(posedge clk_i) begin
         
        if (reset_i) begin
    
          reg_rdata <= #(TCQ) 32'b0;
          reg_rdop <= #(TCQ) 4'b0;
    
         end else begin
    
           case (addr_p1[11:10]) 
             2'b00 : begin
               reg_rdata <= #(TCQ) rdata_t[(32*(0))+31:(32*(0))+0];
               reg_rdop <= #(TCQ) rdop_t[(4*(0))+3:(4*(0))+0];
             end
             2'b01 : begin
               reg_rdata <= #(TCQ) rdata_t[(32*(1))+31:(32*(1))+0];
               reg_rdop <= #(TCQ) rdop_t[(4*(1))+3:(4*(1))+0];
             end
             2'b10 : begin
               reg_rdata <= #(TCQ) rdata_t[(32*(2))+31:(32*(2))+0];
               reg_rdop <= #(TCQ) rdop_t[(4*(2))+3:(4*(2))+0];
             end
             2'b11 : begin
               reg_rdata <= #(TCQ) rdata_t[(32*(3))+31:(32*(3))+0];
               reg_rdop <= #(TCQ) rdop_t[(4*(3))+3:(4*(3))+0];
             end
           endcase
    
          end

        end // always

      end else begin : NOFRMRAMPIPELINE
    
        always @(*) begin

          case (addr_p1[11:10]) 
            2'b00 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(0))+31:(32*(0))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(0))+3:(4*(0))+0];
            end
            2'b01 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(1))+31:(32*(1))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(1))+3:(4*(1))+0];
            end
            2'b10 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(2))+31:(32*(2))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(2))+3:(4*(2))+0];
            end
            2'b11 : begin
              reg_rdata <= #(TCQ) rdata_t[(32*(3))+31:(32*(3))+0];
              reg_rdop <= #(TCQ) rdop_t[(4*(3))+3:(4*(3))+0];
            end
          endcase
    
        end // always

      end // (FROM_RAM_PIPELINE == "TRUE") begin : FRMRAMPIPELINE
  
      assign rdata_o = reg_rdata;
      assign rdop_o = reg_rdop;
      assign baddr = {user_tph_stt_func_num_i[7:0], user_tph_stt_index_i[5:0]};

      always @ (*) begin
    
        if (baddr_p1[13:12] == 2'b00)
          brdata_w = brdata[(32*(0))+31:(32*(0))+0];
        else if (baddr_p1[13:12] == 2'b01)
          brdata_w = brdata[(32*(1))+31:(32*(1))+0];
        else if (baddr_p1[13:12] == 2'b10)
          brdata_w = brdata[(32*(2))+31:(32*(2))+0];
        else
          brdata_w = brdata[(32*(3))+31:(32*(3))+0];
    
      end
    
      assign user_tph_stt_rd_data_o = (baddr_p1[1:0] == 2'b00) ? brdata_w[7:0] : 
                                      (baddr_p1[1:0] == 2'b01) ? brdata_w[15:8] :  
                                      (baddr_p1[1:0] == 2'b10) ? brdata_w[23:16] : brdata_w[31:24];
    
      //
      // BRAM instances
      //

      for (i=0; i<4; i=i+1) begin : BRAM4K

      xp4_usp_smsw_bram_4k_int #(

          .TCQ(TCQ)

        )
        bram_4k_int (
        
          .clk_i (clk_i),
          .reset_i (reset_i),
          .addr_i(addr[9:0]),
          .wdata_i(wdata),
          .wdip_i(wdip),
          .wen_i(bram_4k_wen[(4*i)+3:(4*i)+0]),
          .rdata_o(rdata_t[(32*i)+31:(32*i)+0]),
          .rdop_o(rdop_t[(4*i)+3:(4*i)+0]),
          .baddr_i(baddr[11:2]),
          .brdata_o(brdata[(32*i)+31:(32*i)+0])

        );
        assign bram_4k_wen[(4*i)+3:(4*i)+0] = (i == addr[11:10]) ? wen : 4'h0;
      
      end

    end else begin : TPHR_CAP_NOT_PRESENT 

      assign rdata_o = 32'h0;
      assign rdop_o = 4'h0;
      assign user_tph_stt_rd_data_o = 8'h0;

    end // (PF0_TPHR_CAP_ENABLE == "TRUE") begin : TPHR_CAP_PRESENT

  endgenerate

endmodule
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_512b_intfc.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_512b_intfc #(
     parameter           TCQ = 100
   , parameter           IMPL_TARGET = "SOFT"
   , parameter           AXISTEN_IF_EXT_512_INTFC_RAM_STYLE = "BRAM"
   , parameter           AXISTEN_IF_RQ_CC_REGISTERED_TREADY = "TRUE"
   , parameter           AXI4_USER_DATA_WIDTH = 512
   , parameter           AXI4_CORE_DATA_WIDTH = 256
   , parameter           AXI4_USER_CQ_TUSER_WIDTH = 183
   , parameter           AXI4_USER_CC_TUSER_WIDTH = 81
   , parameter           AXI4_USER_RQ_TUSER_WIDTH = 137
   , parameter           AXI4_USER_RC_TUSER_WIDTH = 161
   , parameter           AXI4_CORE_CQ_TUSER_WIDTH = 88
   , parameter           AXI4_CORE_CC_TUSER_WIDTH = 33
   , parameter           AXI4_CORE_RQ_TUSER_WIDTH = 62
   , parameter           AXI4_CORE_RC_TUSER_WIDTH = 75
   , parameter           AXI4_USER_CQ_TKEEP_WIDTH = 16
   , parameter           AXI4_USER_CC_TKEEP_WIDTH = 16
   , parameter           AXI4_USER_RQ_TKEEP_WIDTH = 16
   , parameter           AXI4_USER_RC_TKEEP_WIDTH = 16
   , parameter           AXI4_CORE_CQ_TKEEP_WIDTH = 8
   , parameter           AXI4_CORE_CC_TKEEP_WIDTH = 8
   , parameter           AXI4_CORE_RQ_TKEEP_WIDTH = 8
   , parameter           AXI4_CORE_RC_TKEEP_WIDTH = 8
   , parameter           AXI4_CORE_CQ_TREADY_WIDTH = 22  
   , parameter           AXI4_CORE_RC_TREADY_WIDTH = 22  
   , parameter           AXISTEN_IF_EXT_512_CQ_STRADDLE="FALSE"
   , parameter           AXISTEN_IF_EXT_512_CC_STRADDLE="FALSE"
   , parameter           AXISTEN_IF_EXT_512_RQ_STRADDLE="FALSE"
   , parameter           AXISTEN_IF_EXT_512_RC_STRADDLE="FALSE"
   , parameter           AXISTEN_IF_EXT_512_RC_4TLP_STRADDLE="TRUE"
   , parameter [1:0]     AXISTEN_IF_CQ_ALIGNMENT_MODE=2'b00
   , parameter [1:0]     AXISTEN_IF_CC_ALIGNMENT_MODE=2'b00
   , parameter [1:0]     AXISTEN_IF_RQ_ALIGNMENT_MODE=2'b00
   , parameter [1:0]     AXISTEN_IF_RC_ALIGNMENT_MODE=2'b00
   , parameter           AXISTEN_IF_RX_PARITY_EN="TRUE"
   , parameter           AXISTEN_IF_TX_PARITY_EN="TRUE"
   ) 
  (
    input  wire           user_clk2_i // 500 MHz clock for core-facing interfaces
   ,input  wire           user_clk_i // 250 MHz clock for client-facing interfaces
   ,input  wire           user_clk_en_i // User clock enable for clock domain crossing
   ,input  wire           reset_n_user_clk_i // Reset in the user clock domain
   ,input  wire           reset_n_user_clk2_i // Reset in the user clock2 domain
   ,input  wire           link_down_reset_i // Link went down
   //-----------------------------------------------------------------------------------------------
   // Client-side interfaces
   //-----------------------------------------------------------------------------------------------
   // CQ Interface
   ,output wire [511:0]   m_axis_cq_tdata_o
   ,output wire           m_axis_cq_tvalid_o
   ,output wire [182:0]   m_axis_cq_tuser_o
   ,output wire           m_axis_cq_tlast_o
   ,output wire [15:0]    m_axis_cq_tkeep_o
   ,input  wire           m_axis_cq_tready_i
   ,input  wire [1:0]     pcie_cq_np_req_i // Client request to deliver NP TLP
   ,output wire [5:0]      pcie_cq_np_req_count_o // Current value of interface credit count for NP TLPs
   // CC Interface
   ,input wire [511:0]    s_axis_cc_tdata_i
   ,input wire            s_axis_cc_tvalid_i
   ,input wire [80:0]     s_axis_cc_tuser_i
   ,input wire            s_axis_cc_tlast_i
   ,input wire [15:0]     s_axis_cc_tkeep_i
   ,output wire            s_axis_cc_tready_o   
   // RQ Interface
   ,input wire [511:0]    s_axis_rq_tdata_i
   ,input wire            s_axis_rq_tvalid_i
   ,input wire [136:0]    s_axis_rq_tuser_i
   ,input wire            s_axis_rq_tlast_i
   ,input wire [15:0]     s_axis_rq_tkeep_i
   ,output wire            s_axis_rq_tready_o   
   // RC Interface
   ,output wire [511:0]   m_axis_rc_tdata_o
   ,output wire           m_axis_rc_tvalid_o
   ,output wire [160:0]   m_axis_rc_tuser_o
   ,output wire           m_axis_rc_tlast_o
   ,output wire [15:0]    m_axis_rc_tkeep_o
   ,input  wire           m_axis_rc_tready_i
   //-----------------------------------------------------------------------------------------------
   // Core-side interfaces
   //-----------------------------------------------------------------------------------------------
   // CQ Interface
   ,input  wire [255:0]   core_cq_tdata_i
   ,input  wire           core_cq_tvalid_i
   ,input  wire [87:0]    core_cq_tuser_i
   ,input  wire           core_cq_tlast_i
   ,input  wire [7:0]     core_cq_tkeep_i
   ,output wire [21:0]     core_cq_tready_o
   ,output wire            posted_req_delivered_o // Signals the delivery of a Posted Req on the CQ interface
   ,output wire            cq_pipeline_empty_o // Indicates that the entire CQ pipeline of the bridge is empty.
   ,output wire            cq_np_user_credit_rcvd_o // Indicates that the user issued one NP credit
   // CC Interface
   ,output wire [255:0]    core_cc_tdata_o
   ,output wire            core_cc_tvalid_o
   ,output wire [32:0]     core_cc_tuser_o
   ,output wire            core_cc_tlast_o
   ,output wire [7:0]      core_cc_tkeep_o
   ,input wire [3:0]      core_cc_tready_i
   // RQ Interface
   ,output wire [255:0]    core_rq_tdata_o
   ,output wire            core_rq_tvalid_o
   ,output wire [61:0]     core_rq_tuser_o
   ,output wire            core_rq_tlast_o
   ,output wire [7:0]      core_rq_tkeep_o
   ,input wire [3:0]      core_rq_tready_i
   // RC Interface
   ,input  wire [255:0]   core_rc_tdata_i
   ,input  wire           core_rc_tvalid_i
   ,input  wire [74:0]    core_rc_tuser_i
   ,input  wire           core_rc_tlast_i
   ,input  wire [7:0]     core_rc_tkeep_i
   ,output wire [21:0]     core_rc_tready_o
   // Completion delivered indications
   ,output wire [1:0]      compl_delivered_o // Completions delivered to user
                                            // 00 = No Compl, 01 = 1 Compl, 11 = 2 Completions
   ,output wire [7:0]      compl_delivered_tag0_o// Tag associated with first delivered Completion
   ,output wire [7:0]      compl_delivered_tag1_o// Tag associated with second delivered Completion
   );

  wire        attr_axisten_if_ext_512_cq_straddle;
  wire        attr_axisten_if_ext_512_cc_straddle;
  wire        attr_axisten_if_ext_512_rq_straddle;
  wire        attr_axisten_if_ext_512_rc_straddle;
  wire        attr_axisten_if_ext_512_rc_4tlp_straddle;
  wire [1:0] attr_axisten_if_cq_alignment_mode;
  wire [1:0] attr_axisten_if_cc_alignment_mode;
  wire [1:0] attr_axisten_if_rq_alignment_mode;
  wire [1:0] attr_axisten_if_rc_alignment_mode;
  wire     attr_axisten_if_rq_cc_registered_tready;
  wire        spare_bit0;
  
  generate
    if (AXISTEN_IF_EXT_512_CQ_STRADDLE == "TRUE")
      assign attr_axisten_if_ext_512_cq_straddle = 1'b1;
    else
      assign attr_axisten_if_ext_512_cq_straddle = 1'b0;
  endgenerate
  
  generate
    if (AXISTEN_IF_EXT_512_CC_STRADDLE == "TRUE")
      assign attr_axisten_if_ext_512_cc_straddle = 1'b1;
    else
      assign attr_axisten_if_ext_512_cc_straddle = 1'b0;
  endgenerate

  generate
    if (AXISTEN_IF_EXT_512_RQ_STRADDLE == "TRUE")
      assign attr_axisten_if_ext_512_rq_straddle = 1'b1;
    else
      assign attr_axisten_if_ext_512_rq_straddle = 1'b0;
  endgenerate

  generate
    if (AXISTEN_IF_EXT_512_RC_STRADDLE == "TRUE")
      assign attr_axisten_if_ext_512_rc_straddle = 1'b1;
    else
      assign attr_axisten_if_ext_512_rc_straddle = 1'b0;
  endgenerate

  generate
    if (AXISTEN_IF_EXT_512_RC_4TLP_STRADDLE == "TRUE")
      assign attr_axisten_if_ext_512_rc_4tlp_straddle = 1'b1;
    else
      assign attr_axisten_if_ext_512_rc_4tlp_straddle = 1'b0;
  endgenerate

  generate
    if (AXISTEN_IF_RQ_CC_REGISTERED_TREADY == "TRUE")
      assign spare_bit0 = 1'b1; 
    else
      assign spare_bit0 = 1'b0; 
  endgenerate
  assign     attr_axisten_if_rq_cc_registered_tready = spare_bit0;

  assign     attr_axisten_if_cq_alignment_mode = AXISTEN_IF_CQ_ALIGNMENT_MODE;
  assign     attr_axisten_if_cc_alignment_mode = AXISTEN_IF_CC_ALIGNMENT_MODE;
  assign     attr_axisten_if_rq_alignment_mode = AXISTEN_IF_RQ_ALIGNMENT_MODE;
  assign     attr_axisten_if_rc_alignment_mode = AXISTEN_IF_RC_ALIGNMENT_MODE;

  xp4_usp_smsw_512b_intfc_int #
    (
     .TCQ(TCQ),
     .IMPL_TARGET(IMPL_TARGET),
     .AXISTEN_IF_EXT_512_INTFC_RAM_STYLE("SRL"),
     .AXI4_USER_DATA_WIDTH(AXI4_USER_DATA_WIDTH),
     .AXI4_CORE_DATA_WIDTH(AXI4_CORE_DATA_WIDTH),
     .AXI4_USER_CQ_TUSER_WIDTH(AXI4_USER_CQ_TUSER_WIDTH),
     .AXI4_USER_CC_TUSER_WIDTH(AXI4_USER_CC_TUSER_WIDTH),
     .AXI4_USER_RQ_TUSER_WIDTH(AXI4_USER_RQ_TUSER_WIDTH),
     .AXI4_USER_RC_TUSER_WIDTH(AXI4_USER_RC_TUSER_WIDTH),
     .AXI4_CORE_CQ_TUSER_WIDTH(AXI4_CORE_CQ_TUSER_WIDTH),
     .AXI4_CORE_CC_TUSER_WIDTH(AXI4_CORE_CC_TUSER_WIDTH),
     .AXI4_CORE_RQ_TUSER_WIDTH(AXI4_CORE_RQ_TUSER_WIDTH),
     .AXI4_CORE_RC_TUSER_WIDTH(AXI4_CORE_RC_TUSER_WIDTH),
     .AXI4_USER_CQ_TKEEP_WIDTH(AXI4_USER_CQ_TKEEP_WIDTH),
     .AXI4_USER_CC_TKEEP_WIDTH(AXI4_USER_CC_TKEEP_WIDTH),
     .AXI4_USER_RQ_TKEEP_WIDTH(AXI4_USER_RQ_TKEEP_WIDTH),
     .AXI4_USER_RC_TKEEP_WIDTH(AXI4_USER_RC_TKEEP_WIDTH),
     .AXI4_CORE_CQ_TKEEP_WIDTH(AXI4_CORE_CQ_TKEEP_WIDTH),
     .AXI4_CORE_CC_TKEEP_WIDTH(AXI4_CORE_CC_TKEEP_WIDTH),
     .AXI4_CORE_RQ_TKEEP_WIDTH(AXI4_CORE_RQ_TKEEP_WIDTH),
     .AXI4_CORE_RC_TKEEP_WIDTH(AXI4_CORE_RC_TKEEP_WIDTH),
     .AXI4_CORE_CQ_TREADY_WIDTH(AXI4_CORE_CQ_TREADY_WIDTH),
     .AXI4_CORE_RC_TREADY_WIDTH(AXI4_CORE_RC_TREADY_WIDTH),
     .AXISTEN_IF_RX_PARITY_EN(AXISTEN_IF_RX_PARITY_EN),
     .AXISTEN_IF_TX_PARITY_EN(AXISTEN_IF_TX_PARITY_EN)
     )
    pcie_4_0_512b_intfc_int_mod
  (
   .user_clk_i         (user_clk_i),
   .user_clk2_i        (user_clk2_i),
   .user_clk_en_i      (user_clk_en_i),
   .reset_n_user_clk_i (reset_n_user_clk_i),
   .reset_n_user_clk2_i(reset_n_user_clk2_i),
   .link_down_reset_i  (link_down_reset_i),
   // Attributes
   .attr_axisten_if_ext_512_cq_straddle_i(attr_axisten_if_ext_512_cq_straddle),
   .attr_axisten_if_ext_512_cc_straddle_i(attr_axisten_if_ext_512_cc_straddle),
   .attr_axisten_if_ext_512_rq_straddle_i(attr_axisten_if_ext_512_rq_straddle),
   .attr_axisten_if_ext_512_rc_straddle_i(attr_axisten_if_ext_512_rc_straddle),
   .attr_axisten_if_ext_512_rc_4tlp_straddle_i(attr_axisten_if_ext_512_rc_4tlp_straddle),
   .attr_axisten_if_cq_alignment_mode_i(attr_axisten_if_cq_alignment_mode),
   .attr_axisten_if_cc_alignment_mode_i(attr_axisten_if_cc_alignment_mode),
   .attr_axisten_if_rq_alignment_mode_i(attr_axisten_if_rq_alignment_mode),
   .attr_axisten_if_rc_alignment_mode_i(attr_axisten_if_rc_alignment_mode),
   .attr_axisten_if_rq_cc_registered_tready_i(attr_axisten_if_rq_cc_registered_tready),
   //-----------------------------------
   // Client-side signals
   //-----------------------------------
   // CQ Interface
   .m_axis_cq_tdata_o  (m_axis_cq_tdata_o),
   .m_axis_cq_tvalid_o (m_axis_cq_tvalid_o),
   .m_axis_cq_tuser_o  (m_axis_cq_tuser_o),
   .m_axis_cq_tlast_o  (m_axis_cq_tlast_o),
   .m_axis_cq_tkeep_o  (m_axis_cq_tkeep_o),
   .m_axis_cq_tready_i (m_axis_cq_tready_i),
   .pcie_cq_np_req_i   (pcie_cq_np_req_i),
   .pcie_cq_np_req_count_o(pcie_cq_np_req_count_o),
   // CC Interface
   .s_axis_cc_tdata_i  (s_axis_cc_tdata_i),
   .s_axis_cc_tvalid_i (s_axis_cc_tvalid_i),
   .s_axis_cc_tuser_i  (s_axis_cc_tuser_i),
   .s_axis_cc_tlast_i  (s_axis_cc_tlast_i),
   .s_axis_cc_tkeep_i  (s_axis_cc_tkeep_i),
   .s_axis_cc_tready_o (s_axis_cc_tready_o),
   // RQ Interface
   .s_axis_rq_tdata_i  (s_axis_rq_tdata_i),
   .s_axis_rq_tvalid_i (s_axis_rq_tvalid_i),
   .s_axis_rq_tuser_i  (s_axis_rq_tuser_i),
   .s_axis_rq_tlast_i  (s_axis_rq_tlast_i),
   .s_axis_rq_tkeep_i  (s_axis_rq_tkeep_i),
   .s_axis_rq_tready_o (s_axis_rq_tready_o),
   // RC Interface
   .m_axis_rc_tdata_o  (m_axis_rc_tdata_o),
   .m_axis_rc_tvalid_o (m_axis_rc_tvalid_o),
   .m_axis_rc_tuser_o  (m_axis_rc_tuser_o),
   .m_axis_rc_tlast_o  (m_axis_rc_tlast_o),
   .m_axis_rc_tkeep_o  (m_axis_rc_tkeep_o),
   .m_axis_rc_tready_i (m_axis_rc_tready_i),
   //-----------------------------------
   // Core-side signals
   //-----------------------------------
   // CQ Interface
   .core_cq_tdata_i    (core_cq_tdata_i),
   .core_cq_tvalid_i   (core_cq_tvalid_i),
   .core_cq_tuser_i    (core_cq_tuser_i),
   .core_cq_tlast_i    (core_cq_tlast_i),
   .core_cq_tkeep_i    (core_cq_tkeep_i),
   .core_cq_tready_o   (core_cq_tready_o),
   .posted_req_delivered_o(posted_req_delivered_o),
   .cq_pipeline_empty_o(cq_pipeline_empty_o),
   .cq_np_user_credit_rcvd_o(cq_np_user_credit_rcvd_o),
   // CC Interface
   .core_cc_tdata_o    (core_cc_tdata_o),
   .core_cc_tvalid_o   (core_cc_tvalid_o),
   .core_cc_tuser_o    (core_cc_tuser_o),
   .core_cc_tlast_o    (core_cc_tlast_o),
   .core_cc_tkeep_o    (core_cc_tkeep_o),
   .core_cc_tready_i   (core_cc_tready_i),
   // RQ Interface
   .core_rq_tdata_o    (core_rq_tdata_o),
   .core_rq_tvalid_o   (core_rq_tvalid_o),
   .core_rq_tuser_o    (core_rq_tuser_o),
   .core_rq_tlast_o    (core_rq_tlast_o),
   .core_rq_tkeep_o    (core_rq_tkeep_o),
   .core_rq_tready_i   (core_rq_tready_i),
   // RC Interface
   .core_rc_tdata_i    (core_rc_tdata_i),
   .core_rc_tvalid_i   (core_rc_tvalid_i),
   .core_rc_tuser_i    (core_rc_tuser_i),
   .core_rc_tlast_i    (core_rc_tlast_i),
   .core_rc_tkeep_i    (core_rc_tkeep_i),
   .core_rc_tready_o   (core_rc_tready_o),
   .compl_delivered_o  (compl_delivered_o),
   .compl_delivered_tag0_o(compl_delivered_tag0_o),
   .compl_delivered_tag1_o(compl_delivered_tag1_o)
   );
endmodule // pcie_4_0_512b_intfc
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_512b_intfc_int.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_512b_intfc_int #(
   parameter TCQ = 100,
   parameter IMPL_TARGET = "SOFT",
   parameter AXISTEN_IF_EXT_512_INTFC_RAM_STYLE = "BRAM",
   parameter AXI4_USER_DATA_WIDTH = 512,
   parameter AXI4_CORE_DATA_WIDTH = 256,
   parameter AXI4_USER_CQ_TUSER_WIDTH = 183,
   parameter AXI4_USER_CC_TUSER_WIDTH = 81,
   parameter AXI4_USER_RQ_TUSER_WIDTH = 137,
   parameter AXI4_USER_RC_TUSER_WIDTH = 161,
   parameter AXI4_CORE_CQ_TUSER_WIDTH = 88,
   parameter AXI4_CORE_CC_TUSER_WIDTH = 33,
   parameter AXI4_CORE_RQ_TUSER_WIDTH = 62,
   parameter AXI4_CORE_RC_TUSER_WIDTH = 75,
   parameter AXI4_USER_CQ_TKEEP_WIDTH = 16,
   parameter AXI4_USER_CC_TKEEP_WIDTH = 16,
   parameter AXI4_USER_RQ_TKEEP_WIDTH = 16,
   parameter AXI4_USER_RC_TKEEP_WIDTH = 16,
   parameter AXI4_CORE_CQ_TKEEP_WIDTH = 8,
   parameter AXI4_CORE_CC_TKEEP_WIDTH = 8,
   parameter AXI4_CORE_RQ_TKEEP_WIDTH = 8,
   parameter AXI4_CORE_RC_TKEEP_WIDTH = 8,
   parameter AXI4_CORE_CQ_TREADY_WIDTH = 22,   
   parameter AXI4_CORE_RC_TREADY_WIDTH = 22,
   parameter AXISTEN_IF_RX_PARITY_EN="TRUE",
   parameter AXISTEN_IF_TX_PARITY_EN="TRUE"
   ) 
  (
    input  wire           user_clk2_i // 500 MHz clock for core-facing interfaces
   ,input  wire           user_clk_i // 250 MHz clock for client-facing interfaces
   ,input  wire           user_clk_en_i // User clock enable for clock domain crossing
   ,input  wire           reset_n_user_clk_i // Reset in the user clock domain
   ,input  wire           reset_n_user_clk2_i // Reset in the user clock2 domain
   ,input  wire           link_down_reset_i // Link went down
   // Attributes
   ,input wire            attr_axisten_if_ext_512_cq_straddle_i // Enable straddle on CQ interface
   ,input wire            attr_axisten_if_ext_512_cc_straddle_i // Enable straddle on CC interface
   ,input wire            attr_axisten_if_ext_512_rq_straddle_i // Enable straddle on RQ interface
   ,input wire            attr_axisten_if_ext_512_rc_straddle_i // Enable straddle on RC interface
   ,input wire            attr_axisten_if_ext_512_rc_4tlp_straddle_i // Enable 4-TLP straddle on RC interface
   ,input wire [1:0]      attr_axisten_if_cq_alignment_mode_i // Alignment mode on CQ interface 
                                                            // (00= Dword-aligned, 10 = 128b address-aligned)
   ,input wire [1:0]      attr_axisten_if_cc_alignment_mode_i // Alignment mode on CC interface 
                                                            // (00 = Dword-aligned, 10 = 128b address-aligned)
   ,input wire [1:0]      attr_axisten_if_rq_alignment_mode_i // Alignment mode on RQ interface 
                                                            // (00 = Dword-aligned, 10 = 128b address-aligned)
   ,input wire [1:0]      attr_axisten_if_rc_alignment_mode_i // Alignment mode on RC interface 
                                                            // (00= Dword-aligned, 10 = 128b address-aligned)
   ,input wire            attr_axisten_if_rq_cc_registered_tready_i // 0 = registered_tready enabled, 1 = registered_tready disabled

   //-----------------------------------------------------------------------------------------------
   // Client-side interfaces
   //-----------------------------------------------------------------------------------------------
   // CQ Interface
   ,output wire [511:0]   m_axis_cq_tdata_o
   ,output wire           m_axis_cq_tvalid_o
   ,output wire [182:0]   m_axis_cq_tuser_o
   ,output wire           m_axis_cq_tlast_o
   ,output wire [15:0]    m_axis_cq_tkeep_o
   ,input  wire           m_axis_cq_tready_i
   ,input  wire [1:0]     pcie_cq_np_req_i // Client request to deliver NP TLP
   ,output wire [5:0]      pcie_cq_np_req_count_o // Current value of interface credit count for NP TLPs
   // CC Interface
   ,input wire [511:0]    s_axis_cc_tdata_i
   ,input wire            s_axis_cc_tvalid_i
   ,input wire [80:0]     s_axis_cc_tuser_i
   ,input wire            s_axis_cc_tlast_i
   ,input wire [15:0]     s_axis_cc_tkeep_i
   ,output wire            s_axis_cc_tready_o   
   // RQ Interface
   ,input wire [511:0]    s_axis_rq_tdata_i
   ,input wire            s_axis_rq_tvalid_i
   ,input wire [136:0]    s_axis_rq_tuser_i
   ,input wire            s_axis_rq_tlast_i
   ,input wire [15:0]     s_axis_rq_tkeep_i
   ,output wire            s_axis_rq_tready_o   
   // RC Interface
   ,output wire [511:0]   m_axis_rc_tdata_o
   ,output wire           m_axis_rc_tvalid_o
   ,output wire [160:0]   m_axis_rc_tuser_o
   ,output wire           m_axis_rc_tlast_o
   ,output wire [15:0]    m_axis_rc_tkeep_o
   ,input  wire           m_axis_rc_tready_i
   //-----------------------------------------------------------------------------------------------
   // Core-side interfaces
   //-----------------------------------------------------------------------------------------------
   // CQ Interface
   ,input  wire [255:0]   core_cq_tdata_i
   ,input  wire           core_cq_tvalid_i
   ,input  wire [87:0]    core_cq_tuser_i
   ,input  wire           core_cq_tlast_i
   ,input  wire [7:0]     core_cq_tkeep_i
   ,output wire [21:0]     core_cq_tready_o
   ,output wire            posted_req_delivered_o // Signals the delivery of a Posted Req on the CQ interface
   ,output wire            cq_pipeline_empty_o // Indicates that the entire CQ pipeline of the bridge is empty.
   ,output wire            cq_np_user_credit_rcvd_o // Indicates that the user issued one NP credit
   // CC Interface
   ,output wire [255:0]    core_cc_tdata_o
   ,output wire            core_cc_tvalid_o
   ,output wire [32:0]     core_cc_tuser_o
   ,output wire            core_cc_tlast_o
   ,output wire [7:0]      core_cc_tkeep_o
   ,input wire [3:0]       core_cc_tready_i
   // RQ Interface
   ,output wire [255:0]    core_rq_tdata_o
   ,output wire            core_rq_tvalid_o
   ,output wire [61:0]     core_rq_tuser_o
   ,output wire            core_rq_tlast_o
   ,output wire [7:0]      core_rq_tkeep_o
   ,input wire [3:0]       core_rq_tready_i
   // RC Interface
   ,input  wire [255:0]   core_rc_tdata_i
   ,input  wire           core_rc_tvalid_i
   ,input  wire [74:0]    core_rc_tuser_i
   ,input  wire           core_rc_tlast_i
   ,input  wire [7:0]     core_rc_tkeep_i
   ,output wire [21:0]     core_rc_tready_o
   // Completion delivered indications
   ,output wire [1:0]      compl_delivered_o // Completions delivered to user
                                            // 00 = No Compl, 01 = 1 Compl, 11 = 2 Completions
   ,output wire [7:0]      compl_delivered_tag0_o// Tag associated with first delivered Completion
   ,output wire [7:0]      compl_delivered_tag1_o// Tag associated with second delivered Completion
   );

  // CQ Module
  xp4_usp_smsw_512b_cq_intfc #
    (
     .TCQ(TCQ),
     .IMPL_TARGET(IMPL_TARGET),
     .AXISTEN_IF_EXT_512_INTFC_RAM_STYLE(AXISTEN_IF_EXT_512_INTFC_RAM_STYLE),
     .AXI4_USER_DATA_WIDTH(AXI4_USER_DATA_WIDTH),
     .AXI4_CORE_DATA_WIDTH(AXI4_CORE_DATA_WIDTH),
     .AXI4_USER_CQ_TUSER_WIDTH(AXI4_USER_CQ_TUSER_WIDTH),
     .AXI4_CORE_CQ_TUSER_WIDTH(AXI4_CORE_CQ_TUSER_WIDTH),
     .AXI4_USER_CQ_TKEEP_WIDTH(AXI4_USER_CQ_TKEEP_WIDTH),
     .AXI4_CORE_CQ_TKEEP_WIDTH(AXI4_CORE_CQ_TKEEP_WIDTH),
     .AXI4_CORE_CQ_TREADY_WIDTH(AXI4_CORE_CQ_TREADY_WIDTH),
     .PARITY_ENABLE(1)
     ) 
    pcie_4_0_512b_cq_intfc_mod
   (
    .user_clk2_i        (user_clk2_i),
    .user_clk_i         (user_clk_i),
    .user_clk_en_i      (user_clk_en_i),
    .reset_n_user_clk_i (reset_n_user_clk_i),
    .reset_n_user_clk2_i(reset_n_user_clk2_i),
    .link_down_reset_i  (link_down_reset_i),
   // Attributes
    .attr_straddle_en_i (attr_axisten_if_ext_512_cq_straddle_i),
    .attr_alignment_mode_i(attr_axisten_if_cq_alignment_mode_i),
   //-----------------------------------------------------------------------------------------------
   // Client-side signals
   //-----------------------------------------------------------------------------------------------
    .m_axis_cq_tdata_o  (m_axis_cq_tdata_o),
    .m_axis_cq_tvalid_o (m_axis_cq_tvalid_o),
    .m_axis_cq_tuser_o  (m_axis_cq_tuser_o),
    .m_axis_cq_tlast_o  (m_axis_cq_tlast_o),
    .m_axis_cq_tkeep_o  (m_axis_cq_tkeep_o),
    .m_axis_cq_tready_i (m_axis_cq_tready_i),
    .pcie_cq_np_req_i   (pcie_cq_np_req_i), 
    .pcie_cq_np_req_count_o(pcie_cq_np_req_count_o),
   //-----------------------------------------------------------------------------------------------
   // Core-side signals
   //-----------------------------------------------------------------------------------------------
    .core_cq_tdata_i    (core_cq_tdata_i),
    .core_cq_tvalid_i   (core_cq_tvalid_i),
    .core_cq_tuser_i    (core_cq_tuser_i),
    .core_cq_tlast_i    (core_cq_tlast_i),
    .core_cq_tkeep_i    (core_cq_tkeep_i),
    .core_cq_tready_o   (core_cq_tready_o),
    .posted_req_delivered_o(posted_req_delivered_o),
    .cq_pipeline_empty_o(cq_pipeline_empty_o),
    .cq_np_user_credit_rcvd_o(cq_np_user_credit_rcvd_o)
    );
  
  // CC Module
  xp4_usp_smsw_512b_cc_intfc #
    (
     .TCQ(TCQ),
     .IMPL_TARGET(IMPL_TARGET),
     .AXI4_USER_DATA_WIDTH(AXI4_USER_DATA_WIDTH),
     .AXI4_CORE_DATA_WIDTH(AXI4_CORE_DATA_WIDTH),
     .AXI4_USER_CC_TUSER_WIDTH(AXI4_USER_CC_TUSER_WIDTH),
     .AXI4_CORE_CC_TUSER_WIDTH(AXI4_CORE_CC_TUSER_WIDTH),
     .AXI4_USER_CC_TKEEP_WIDTH(AXI4_USER_CC_TKEEP_WIDTH),
     .AXI4_CORE_CC_TKEEP_WIDTH(AXI4_CORE_CC_TKEEP_WIDTH),
     .PARITY_ENABLE(1)
     ) 
    pcie_4_0_512b_cc_intfc_mod
   (
    .user_clk2_i        (user_clk2_i),
    .user_clk_i         (user_clk_i),
    .user_clk_en_i      (user_clk_en_i),
    .reset_n_user_clk_i (reset_n_user_clk_i),
    .reset_n_user_clk2_i(reset_n_user_clk2_i),
    .link_down_reset_i  (link_down_reset_i),
   // Attributes
    .attr_straddle_en_i (attr_axisten_if_ext_512_cc_straddle_i),
    .attr_alignment_mode_i(attr_axisten_if_cc_alignment_mode_i),
    .attr_axisten_if_rq_cc_registered_tready_i(attr_axisten_if_rq_cc_registered_tready_i),
   //-----------------------------------------------------------------------------------------------
   // Client-side signals
   //-----------------------------------------------------------------------------------------------
    .s_axis_cc_tdata_i  (s_axis_cc_tdata_i),
    .s_axis_cc_tvalid_i (s_axis_cc_tvalid_i),
    .s_axis_cc_tuser_i  (s_axis_cc_tuser_i),
    .s_axis_cc_tlast_i  (s_axis_cc_tlast_i),
    .s_axis_cc_tkeep_i  (s_axis_cc_tkeep_i),
    .s_axis_cc_tready_o (s_axis_cc_tready_o),   
   //-----------------------------------------------------------------------------------------------
   // Core-side signals
   //-----------------------------------------------------------------------------------------------
    .core_cc_tdata_o  (core_cc_tdata_o),
    .core_cc_tvalid_o (core_cc_tvalid_o),
    .core_cc_tuser_o  (core_cc_tuser_o),
    .core_cc_tlast_o  (core_cc_tlast_o),
    .core_cc_tkeep_o  (core_cc_tkeep_o),
    .core_cc_tready_i (core_cc_tready_i)
    );

  // RQ Module
  xp4_usp_smsw_512b_rq_intfc #
    (
     .TCQ(TCQ),
     .IMPL_TARGET(IMPL_TARGET),
     .AXI4_USER_DATA_WIDTH(AXI4_USER_DATA_WIDTH),
     .AXI4_CORE_DATA_WIDTH(AXI4_CORE_DATA_WIDTH),
     .AXI4_USER_RQ_TUSER_WIDTH(AXI4_USER_RQ_TUSER_WIDTH),
     .AXI4_CORE_RQ_TUSER_WIDTH(AXI4_CORE_RQ_TUSER_WIDTH),
     .AXI4_USER_RQ_TKEEP_WIDTH(AXI4_USER_RQ_TKEEP_WIDTH),
     .AXI4_CORE_RQ_TKEEP_WIDTH(AXI4_CORE_RQ_TKEEP_WIDTH),
     .PARITY_ENABLE(1)
     ) 
    pcie_4_0_512b_rq_intfc_mod
   (
    .user_clk2_i        (user_clk2_i),
    .user_clk_i         (user_clk_i),
    .user_clk_en_i      (user_clk_en_i),
    .reset_n_user_clk_i (reset_n_user_clk_i),
    .reset_n_user_clk2_i(reset_n_user_clk2_i),
    .link_down_reset_i  (link_down_reset_i),
   // Attributes
    .attr_straddle_en_i (attr_axisten_if_ext_512_rq_straddle_i),
    .attr_alignment_mode_i(attr_axisten_if_rq_alignment_mode_i),
    .attr_axisten_if_rq_cc_registered_tready_i(attr_axisten_if_rq_cc_registered_tready_i),
   //-----------------------------------------------------------------------------------------------
   // Client-side signals
   //-----------------------------------------------------------------------------------------------
    .s_axis_rq_tdata_i  (s_axis_rq_tdata_i),
    .s_axis_rq_tvalid_i (s_axis_rq_tvalid_i),
    .s_axis_rq_tuser_i  (s_axis_rq_tuser_i),
    .s_axis_rq_tlast_i  (s_axis_rq_tlast_i),
    .s_axis_rq_tkeep_i  (s_axis_rq_tkeep_i),
    .s_axis_rq_tready_o (s_axis_rq_tready_o),   
   //-----------------------------------------------------------------------------------------------
   // Core-side signals
   //-----------------------------------------------------------------------------------------------
    .core_rq_tdata_o  (core_rq_tdata_o),
    .core_rq_tvalid_o (core_rq_tvalid_o),
    .core_rq_tuser_o  (core_rq_tuser_o),
    .core_rq_tlast_o  (core_rq_tlast_o),
    .core_rq_tkeep_o  (core_rq_tkeep_o),
    .core_rq_tready_i  (core_rq_tready_i)
    );

  // RC Module
  xp4_usp_smsw_512b_rc_intfc #
    (
     .TCQ(TCQ),
     .IMPL_TARGET(IMPL_TARGET),
     .AXI4_USER_DATA_WIDTH(AXI4_USER_DATA_WIDTH),
     .AXI4_CORE_DATA_WIDTH(AXI4_CORE_DATA_WIDTH),
     .AXI4_USER_RC_TUSER_WIDTH(AXI4_USER_RC_TUSER_WIDTH),
     .AXI4_CORE_RC_TUSER_WIDTH(AXI4_CORE_RC_TUSER_WIDTH),
     .AXI4_USER_RC_TKEEP_WIDTH(AXI4_USER_RC_TKEEP_WIDTH),
     .AXI4_CORE_RC_TKEEP_WIDTH(AXI4_CORE_RC_TKEEP_WIDTH),
     .AXI4_CORE_RC_TREADY_WIDTH(AXI4_CORE_RC_TREADY_WIDTH),
     .PARITY_ENABLE(1)
     ) 
    pcie_4_0_512b_rc_intfc_mod
   (
    .user_clk2_i        (user_clk2_i),
    .user_clk_i         (user_clk_i),
    .user_clk_en_i      (user_clk_en_i),
    .reset_n_user_clk_i (reset_n_user_clk_i),
    .reset_n_user_clk2_i(reset_n_user_clk2_i),
    .link_down_reset_i  (link_down_reset_i),
   // Attributes
    .attr_straddle_en_i (attr_axisten_if_ext_512_rc_straddle_i),
    .attr_4tlp_straddle_en_i (attr_axisten_if_ext_512_rc_4tlp_straddle_i),
    .attr_alignment_mode_i(attr_axisten_if_rc_alignment_mode_i),
   //-----------------------------------------------------------------------------------------------
   // Client-side signals
   //-----------------------------------------------------------------------------------------------
    .m_axis_rc_tdata_o  (m_axis_rc_tdata_o),
    .m_axis_rc_tvalid_o (m_axis_rc_tvalid_o),
    .m_axis_rc_tuser_o  (m_axis_rc_tuser_o),
    .m_axis_rc_tlast_o  (m_axis_rc_tlast_o),
    .m_axis_rc_tkeep_o  (m_axis_rc_tkeep_o),
    .m_axis_rc_tready_i (m_axis_rc_tready_i),
   //-----------------------------------------------------------------------------------------------
   // Core-side signals
   //-----------------------------------------------------------------------------------------------
    .core_rc_tdata_i    (core_rc_tdata_i),
    .core_rc_tvalid_i   (core_rc_tvalid_i),
    .core_rc_tuser_i    (core_rc_tuser_i),
    .core_rc_tlast_i    (core_rc_tlast_i),
    .core_rc_tkeep_i    (core_rc_tkeep_i),
    .core_rc_tready_o   (core_rc_tready_o),
   // Completion delivered indications
    .compl_delivered_o  (compl_delivered_o),
    .compl_delivered_tag0_o(compl_delivered_tag0_o),
    .compl_delivered_tag1_o(compl_delivered_tag1_o)
    );

endmodule // pcie_4_0_512b_intfc_int
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_512b_async_fifo.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_512b_async_fifo #(
   parameter TCQ = 100,
   parameter IMPL_TARGET = "SOFT",
   parameter IN_DATA_WIDTH = 512,
   parameter FIFO_WIDTH = 256,
   parameter FIFO_DEPTH = 16,
   parameter FIFO_ALMOST_FULL_THRESHOLD = 7
   ) 
  (
   // Write side
    input  wire           clk_i // clock
   ,input  wire           clk_en_i // clock enable, valid in alternate cycles
   ,input  wire           reset_n_i // Reset 
   ,input  wire           link_down_reset_i // Reset FIFO on link down
   ,input wire [IN_DATA_WIDTH-1:0] write_data_i
   ,input wire [1:0]       write_en_i
   ,output wire            fifo_almost_full_o
   // Read side
   ,input                 read_en_i
   ,output wire [FIFO_WIDTH-1:0] read_data_o
   ,output wire           read_data_valid_o
   );
   
  reg [3:0]    read_ptr;
  reg [3:0]    fifo_occupancy;
  reg            fifo_empty;

  integer    i;

  reg [FIFO_WIDTH-1:0]  ram_array[FIFO_DEPTH-1:0];
  reg [FIFO_WIDTH-1:0]     write_data_reg;
  reg             write_data_valid_reg;

  // Convert input data to core clock domain by registering it.
  // Serialize writes of lower and upper halves.
  
  always @(posedge clk_i)
    if (~reset_n_i)
      write_data_reg <= #TCQ {FIFO_WIDTH{1'b0}};
    else
      begin
    if (~clk_en_i & write_en_i[0])
      write_data_reg[FIFO_WIDTH-1:0] <= #TCQ write_data_i[IN_DATA_WIDTH/2-1:0];
    else if (clk_en_i & write_en_i[1])
      write_data_reg[FIFO_WIDTH-1:0] <= #TCQ write_data_i[IN_DATA_WIDTH-1:IN_DATA_WIDTH/2];
      end

  always @(posedge clk_i)
    if (~reset_n_i)
      write_data_valid_reg <= #TCQ 1'b0;
    else
      begin
    if (~clk_en_i)
      write_data_valid_reg <= #TCQ  write_en_i[0];
    else
      write_data_valid_reg <= #TCQ  write_en_i[1];
      end

  // synthesis translate_off
  initial
  begin
    for (i=0; i < FIFO_WIDTH; i=i+1)
      begin
    ram_array[i] = 0;
      end
  end
  // synthesis translate_on

  //Write to SRL inputs, and shift SRL
  always @(posedge clk_i)
    if (write_data_valid_reg)
      begin
    for (i= (FIFO_DEPTH-1); i>0; i=i-1)
      ram_array[i] <= #TCQ ram_array[i-1];
     ram_array[0]   <= #TCQ write_data_reg[FIFO_WIDTH-1:0];
      end
    
   // Read pointer
   always @(posedge clk_i)
     if (~reset_n_i)
       read_ptr <= #(TCQ) 4'd0;
     else if (link_down_reset_i)
       read_ptr <= #(TCQ) 4'd0;
     else if ((read_en_i & ~fifo_empty) &
          (~write_data_valid_reg))
       // Read but no write in this cycle
       begin
     if (read_ptr != 4'd0)
       read_ptr <= #TCQ read_ptr - 4'd1;
       end
       else if (~(read_en_i & ~fifo_empty) &
          write_data_valid_reg)
     // Write but no read in this cycle
     begin
       if (~fifo_empty)
         read_ptr <= #TCQ read_ptr + 4'd1;
     end
  
   // Maintain FIFO occupancy
   always @(posedge clk_i)
     if (~reset_n_i)
       begin
     fifo_occupancy <= #TCQ 4'd0;
     fifo_empty <= #TCQ 1'b1;
       end
     else if (link_down_reset_i)
       begin
     fifo_occupancy <= #TCQ 4'd0;
     fifo_empty <= #TCQ 1'b1;
       end
     else if ((read_en_i & ~fifo_empty) &
          (~write_data_valid_reg))
       // Read but no write in this cycle
       begin
     fifo_occupancy <= #TCQ fifo_occupancy - 4'd1;
     fifo_empty <= #TCQ (fifo_occupancy == 4'd1);
       end
     else if (~(read_en_i & ~fifo_empty) &
          write_data_valid_reg)
       // Write but no read in this cycle
       begin
     fifo_occupancy <= #TCQ fifo_occupancy + 4'd1;
     fifo_empty <= #TCQ 1'b0;
       end
  
  assign fifo_almost_full_o = (fifo_occupancy >= FIFO_ALMOST_FULL_THRESHOLD);

   assign    read_data_o = ram_array[read_ptr[3:0]];
   assign    read_data_valid_o = ~fifo_empty;

endmodule // pcie_4_0_512b_async_fifo




//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_512b_cc_intfc.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_512b_cc_intfc #(
   parameter TCQ = 100,
   parameter IMPL_TARGET = "SOFT",
   parameter AXI4_USER_DATA_WIDTH = 512,
   parameter AXI4_CORE_DATA_WIDTH = 256,
   parameter AXI4_USER_CC_TUSER_WIDTH = 81,
   parameter AXI4_CORE_CC_TUSER_WIDTH = 33,
   parameter AXI4_USER_CC_TKEEP_WIDTH = 16,
   parameter AXI4_CORE_CC_TKEEP_WIDTH = 8,
   parameter AXI4_CORE_CC_TREADY_WIDTH = 4,
   parameter PARITY_ENABLE = 0
   ) 
  (
    input  wire           user_clk2_i // 500 MHz clock for core-facing interfaces
   ,input  wire           user_clk_i // 250 MHz clock for client-facing interfaces
   ,input  wire           user_clk_en_i // User clock enable for clock domain crossing
   ,input  wire           reset_n_user_clk_i // Reset in the user clock domain
   ,input  wire           reset_n_user_clk2_i // Reset in the user clock2 domain
   ,input  wire           link_down_reset_i // Link went down
   // Attributes
   ,input  wire           attr_straddle_en_i // Enable straddle
   ,input wire [1:0]      attr_alignment_mode_i // Payload alignment mode
                                                // (00= Dword-aligned, 10 = 128b address-aligned)
   ,input wire            attr_axisten_if_rq_cc_registered_tready_i // 0 = registered_tready enabled, 1 = registered_tready disabled
   //-----------------------------------------------------------------------------------------------
   // Client-side signals
   //-----------------------------------------------------------------------------------------------
   ,input wire [AXI4_USER_DATA_WIDTH-1:0]    s_axis_cc_tdata_i
   ,input wire            s_axis_cc_tvalid_i
   ,input wire [AXI4_USER_CC_TUSER_WIDTH-1:0]     s_axis_cc_tuser_i
   ,input wire            s_axis_cc_tlast_i
   ,input wire [AXI4_USER_CC_TKEEP_WIDTH-1:0]     s_axis_cc_tkeep_i
   ,output reg            s_axis_cc_tready_o   
   //-----------------------------------------------------------------------------------------------
   // Core-side signals
   //-----------------------------------------------------------------------------------------------
   ,output wire [AXI4_CORE_DATA_WIDTH-1:0]    core_cc_tdata_o
   ,output wire            core_cc_tvalid_o
   ,output wire [AXI4_CORE_CC_TUSER_WIDTH-1:0]   core_cc_tuser_o
   ,output wire            core_cc_tlast_o
   ,output wire [AXI4_CORE_CC_TKEEP_WIDTH-1:0]   core_cc_tkeep_o
   ,input wire [AXI4_CORE_CC_TREADY_WIDTH-1:0] core_cc_tready_i
   );

   localparam FIFO_IN_DATA_WIDTH = AXI4_USER_DATA_WIDTH + AXI4_USER_CC_TKEEP_WIDTH + AXI4_CORE_CC_TUSER_WIDTH*2 +
                   2;
   localparam FIFO_OUT_DATA_WIDTH = FIFO_IN_DATA_WIDTH/2;

   localparam OUTPUT_MUX_IN_DATA_WIDTH = AXI4_CORE_DATA_WIDTH + AXI4_CORE_CC_TKEEP_WIDTH + AXI4_CORE_CC_TUSER_WIDTH + 1;

   reg [AXI4_USER_DATA_WIDTH-1:0] s_axis_cc_tdata_reg;
   reg                   s_axis_cc_tvalid_reg_lower;
   reg                   s_axis_cc_tvalid_reg_upper;
   reg [AXI4_USER_CC_TKEEP_WIDTH-1:0] s_axis_cc_tkeep_reg;
   reg                       s_axis_cc_tlast_reg_lower;
   reg                       s_axis_cc_tlast_reg_upper;
   reg [AXI4_USER_CC_TUSER_WIDTH-1:0] s_axis_cc_tuser_reg;

   wire [1:0]                   s_axis_cc_sop;
   wire [1:0]                   s_axis_cc_eop;
   wire [1:0]                   s_axis_cc_sop0_ptr;
   wire [3:0]                   s_axis_cc_eop0_ptr;
   wire [3:0]                   s_axis_cc_eop1_ptr;
   wire [63:0]                   s_axis_cc_parity;

   wire [AXI4_CORE_CC_TUSER_WIDTH*2-1:0] fifo_in_data_tuser;
   wire [1:0]                  fifo_in_data_tlast;

  wire [FIFO_IN_DATA_WIDTH-1:0]      fifo_in_data;
   wire [1:0]                 fifo_in_data_valid;
   wire                  fifo_almost_full_user_clk;

   reg                      s_axis_cc_tuser_discontinue_reg_lower;
   reg                      s_axis_cc_tuser_discontinue_reg_upper;

  wire [FIFO_OUT_DATA_WIDTH-1:0]      fifo_read_data;
   wire                  fifo_read_data_valid;
   wire                  output_mux_ready;

  reg [AXI4_CORE_CC_TREADY_WIDTH-1:0]      core_cc_tready_reg;
  wire [AXI4_CORE_CC_TREADY_WIDTH-1:0]      core_cc_tready_int;

   // Register input data

  assign                  s_axis_cc_sop[1:0] =  s_axis_cc_tuser_i[1:0];
  assign                  s_axis_cc_sop0_ptr[1:0] =  s_axis_cc_tuser_i[3:2];
  assign                  s_axis_cc_eop[1:0] =  s_axis_cc_tuser_i[7:6];
  assign                  s_axis_cc_eop0_ptr[3:0] =  s_axis_cc_tuser_i[11:8];
  assign                  s_axis_cc_eop1_ptr[3:0] =  s_axis_cc_tuser_i[15:12];

   always @(posedge user_clk_i)
     if (~reset_n_user_clk_i)
       begin
      s_axis_cc_tdata_reg <= {AXI4_USER_DATA_WIDTH{1'b0}};
      s_axis_cc_tvalid_reg_lower <= 1'b0;
      s_axis_cc_tvalid_reg_upper <= 1'b0;
      s_axis_cc_tkeep_reg <= {AXI4_USER_CC_TKEEP_WIDTH{1'b0}};
      s_axis_cc_tuser_reg <= {AXI4_USER_CC_TUSER_WIDTH{1'b0}};
     s_axis_cc_tuser_discontinue_reg_lower <= 1'b0;
     s_axis_cc_tuser_discontinue_reg_upper <= 1'b0;
     s_axis_cc_tlast_reg_lower <= 1'b0;
     s_axis_cc_tlast_reg_upper <= 1'b0;
       end
     else
       begin
      s_axis_cc_tdata_reg <= s_axis_cc_tdata_i;
      s_axis_cc_tvalid_reg_lower <= s_axis_cc_tvalid_i & s_axis_cc_tready_o;
      s_axis_cc_tvalid_reg_upper <= attr_straddle_en_i? s_axis_cc_tvalid_i & s_axis_cc_tready_o &
                    (~s_axis_cc_eop[0] | s_axis_cc_eop0_ptr[3] |
                     (s_axis_cc_sop[0] & s_axis_cc_sop0_ptr[1]) |
                     s_axis_cc_sop[1]):
                    s_axis_cc_tvalid_i & s_axis_cc_tready_o &
                    (~s_axis_cc_tlast_i | s_axis_cc_tkeep_i[8]);
     // Generate tkeep settings for core side
     if (~attr_straddle_en_i)
       s_axis_cc_tkeep_reg[7:0] <= s_axis_cc_tkeep_i[7:0];
     else if (s_axis_cc_tvalid_i & s_axis_cc_tready_o)
       begin
         if (~s_axis_cc_eop[0] | s_axis_cc_eop0_ptr[3])
           s_axis_cc_tkeep_reg[7:0] <= 8'hff;
         else
           case(s_axis_cc_eop0_ptr[2:0])
         3'd0: s_axis_cc_tkeep_reg[7:0] <= 8'h01;
         3'd1: s_axis_cc_tkeep_reg[7:0] <= 8'h03;
         3'd2: s_axis_cc_tkeep_reg[7:0] <= 8'h07;
         3'd3: s_axis_cc_tkeep_reg[7:0] <= 8'h0f;
         3'd4: s_axis_cc_tkeep_reg[7:0] <= 8'h1f;
         3'd5: s_axis_cc_tkeep_reg[7:0] <= 8'h3f;
         3'd6: s_axis_cc_tkeep_reg[7:0] <= 8'h7f;
         default: s_axis_cc_tkeep_reg[7:0] <= 8'hff;
           endcase // case(s_axis_cc_eop0_ptr[2:0])
       end // if (s_axis_cc_tvalid_i & s_axis_cc_tready_o)
     else
       s_axis_cc_tkeep_reg[7:0] <= 8'd0;
         
     if (~attr_straddle_en_i)
       s_axis_cc_tkeep_reg[15:8] <= s_axis_cc_tkeep_i[15:8];
     else if (s_axis_cc_tvalid_i & s_axis_cc_tready_o)
       begin
         if (~s_axis_cc_eop[0])
           s_axis_cc_tkeep_reg[15:8] <= 8'hff;
         else if (s_axis_cc_eop0_ptr[3])
           case(s_axis_cc_eop0_ptr[2:0])
         3'd0: s_axis_cc_tkeep_reg[15:8] <= 8'h01;
         3'd1: s_axis_cc_tkeep_reg[15:8] <= 8'h03;
         3'd2: s_axis_cc_tkeep_reg[15:8] <= 8'h07;
         3'd3: s_axis_cc_tkeep_reg[15:8] <= 8'h0f;
         3'd4: s_axis_cc_tkeep_reg[15:8] <= 8'h1f;
         3'd5: s_axis_cc_tkeep_reg[15:8] <= 8'h3f;
         3'd6: s_axis_cc_tkeep_reg[15:8] <= 8'h7f;
         default: s_axis_cc_tkeep_reg[15:8] <= 8'hff;
           endcase // case(s_axis_cc_eop0_ptr[2:0])
         else if ((s_axis_cc_sop[0] && (s_axis_cc_sop0_ptr[1]))||
              s_axis_cc_sop[1])
           // Packet starting in second half
           begin
         if (~s_axis_cc_eop[1])
           s_axis_cc_tkeep_reg[15:8] <= 8'hff;
         else
           case(s_axis_cc_eop1_ptr[2:0])
             3'd2: s_axis_cc_tkeep_reg[15:8] <= 8'h07;
             3'd3: s_axis_cc_tkeep_reg[15:8] <= 8'h0f;
             3'd4: s_axis_cc_tkeep_reg[15:8] <= 8'h1f;
             3'd5: s_axis_cc_tkeep_reg[15:8] <= 8'h3f;
             3'd6: s_axis_cc_tkeep_reg[15:8] <= 8'h7f;
             default: s_axis_cc_tkeep_reg[15:8] <= 8'hff;
           endcase // case(s_axis_cc_eop1_ptr[2:0])
           end // if ((s_axis_cc_sop[0] && (s_axis_cc_sop0_ptr[1]))||...
         else
           s_axis_cc_tkeep_reg[15:8] <= 8'd0;
       end // if (s_axis_cc_tvalid_i & s_axis_cc_tready_o)
     else
       s_axis_cc_tkeep_reg[15:8] <= 8'd0;

      s_axis_cc_tuser_reg <= s_axis_cc_tuser_i;
     // Generate discontinue for lower and upper halves
     if (~attr_straddle_en_i) 
       begin
         s_axis_cc_tuser_discontinue_reg_lower <= s_axis_cc_tuser_i[16] &
                              (~s_axis_cc_tlast_i |
                               ~s_axis_cc_tkeep_i[8]);
         s_axis_cc_tuser_discontinue_reg_upper <= s_axis_cc_tuser_i[16] &
                              (~s_axis_cc_tlast_i |
                               s_axis_cc_tkeep_i[8]);
       end // if (~attr_straddle_en_i)
     else
       begin
         s_axis_cc_tuser_discontinue_reg_lower <= s_axis_cc_tuser_i[16] &
                              (~s_axis_cc_eop[0] |
                               ~s_axis_cc_eop0_ptr[3]);
         s_axis_cc_tuser_discontinue_reg_upper <= s_axis_cc_tuser_i[16] &
                              (~s_axis_cc_eop[0] |
                               s_axis_cc_eop0_ptr[3]);
       end // else: !if(~attr_straddle_en_i)

     // Generate tlast for lower and upper halves
     s_axis_cc_tlast_reg_lower <= attr_straddle_en_i? (s_axis_cc_eop[0] & ~s_axis_cc_eop0_ptr[3]):
                      s_axis_cc_tlast_i & ~s_axis_cc_tkeep_i[8];
     s_axis_cc_tlast_reg_upper <= attr_straddle_en_i? (s_axis_cc_eop[0] & s_axis_cc_eop0_ptr[3]) |
                      s_axis_cc_eop[1]:
                      s_axis_cc_tlast_i & s_axis_cc_tkeep_i[8];
       end // else: !if(~reset_n_user_clk_i)

  assign  s_axis_cc_parity[63:0] =  PARITY_ENABLE? s_axis_cc_tuser_reg[80:17] : 64'd0;

   // Generate the tuser signals for the core side
   // discontinue
  assign  fifo_in_data_tuser[0] = s_axis_cc_tuser_discontinue_reg_lower;
  assign  fifo_in_data_tuser[AXI4_CORE_CC_TUSER_WIDTH+0] = s_axis_cc_tuser_discontinue_reg_upper;
   // parity
   assign fifo_in_data_tuser[32:1] = s_axis_cc_parity[31:0];
   assign fifo_in_data_tuser[AXI4_CORE_CC_TUSER_WIDTH+32:AXI4_CORE_CC_TUSER_WIDTH+1] = s_axis_cc_parity[63:32];
   
   // Generate tlast for lower and upper halves
  assign fifo_in_data_tlast[0] = s_axis_cc_tlast_reg_lower;
  assign fifo_in_data_tlast[1] = s_axis_cc_tlast_reg_upper;
   
   // Generate valid for upper half
  assign fifo_in_data_valid[0] = s_axis_cc_tvalid_reg_lower;
  assign fifo_in_data_valid[1] = s_axis_cc_tvalid_reg_upper;

   assign fifo_in_data[AXI4_CORE_DATA_WIDTH-1:0] = s_axis_cc_tdata_reg[AXI4_CORE_DATA_WIDTH-1:0];
   assign fifo_in_data[FIFO_IN_DATA_WIDTH/2+AXI4_CORE_DATA_WIDTH-1:FIFO_IN_DATA_WIDTH/2] =
      s_axis_cc_tdata_reg[AXI4_CORE_DATA_WIDTH*2-1:AXI4_CORE_DATA_WIDTH];

   assign fifo_in_data[AXI4_CORE_DATA_WIDTH + AXI4_CORE_CC_TKEEP_WIDTH-1: AXI4_CORE_DATA_WIDTH] =
      s_axis_cc_tkeep_reg[AXI4_CORE_CC_TKEEP_WIDTH-1:0];
  assign  fifo_in_data[FIFO_IN_DATA_WIDTH/2 + AXI4_CORE_DATA_WIDTH + AXI4_CORE_CC_TKEEP_WIDTH-1:
               FIFO_IN_DATA_WIDTH/2 + AXI4_CORE_DATA_WIDTH] =
      s_axis_cc_tkeep_reg[AXI4_CORE_CC_TKEEP_WIDTH*2-1:AXI4_CORE_CC_TKEEP_WIDTH];

   assign fifo_in_data[AXI4_CORE_DATA_WIDTH + AXI4_CORE_CC_TKEEP_WIDTH +  AXI4_CORE_CC_TUSER_WIDTH-1:
               AXI4_CORE_DATA_WIDTH + AXI4_CORE_CC_TKEEP_WIDTH] = 
      fifo_in_data_tuser[AXI4_CORE_CC_TUSER_WIDTH-1:0];
   assign fifo_in_data[FIFO_IN_DATA_WIDTH/2 + AXI4_CORE_DATA_WIDTH + AXI4_CORE_CC_TKEEP_WIDTH +  AXI4_CORE_CC_TUSER_WIDTH-1:
               FIFO_IN_DATA_WIDTH/2 + AXI4_CORE_DATA_WIDTH + AXI4_CORE_CC_TKEEP_WIDTH] = 
      fifo_in_data_tuser[AXI4_CORE_CC_TUSER_WIDTH*2-1:AXI4_CORE_CC_TUSER_WIDTH];

   assign fifo_in_data[AXI4_CORE_DATA_WIDTH + AXI4_CORE_CC_TKEEP_WIDTH +  AXI4_CORE_CC_TUSER_WIDTH] =
      fifo_in_data_tlast[0];
   assign fifo_in_data[FIFO_IN_DATA_WIDTH/2 + AXI4_CORE_DATA_WIDTH + AXI4_CORE_CC_TKEEP_WIDTH +  AXI4_CORE_CC_TUSER_WIDTH] =
      fifo_in_data_tlast[1];

   // De-assert ready when FIFO is almost full
   always @(posedge user_clk_i)
     if (~reset_n_user_clk_i)
       s_axis_cc_tready_o <= 1'b0;
     else
       s_axis_cc_tready_o <= #(TCQ) ~fifo_almost_full_user_clk;

  // Register tready from hard block
   always @(posedge user_clk2_i)
     if (~reset_n_user_clk2_i)
       core_cc_tready_reg <= {AXI4_CORE_CC_TREADY_WIDTH{1'b0}};
     else
       core_cc_tready_reg <= core_cc_tready_i;

  assign  core_cc_tready_int = attr_axisten_if_rq_cc_registered_tready_i?
      core_cc_tready_reg : core_cc_tready_i;

   // Async FIFO
   xp4_usp_smsw_512b_async_fifo #
     (
      .TCQ(TCQ),
      .IMPL_TARGET(IMPL_TARGET),
      .IN_DATA_WIDTH(FIFO_IN_DATA_WIDTH),
      .FIFO_WIDTH(FIFO_OUT_DATA_WIDTH),
      .FIFO_DEPTH(16),
      .FIFO_ALMOST_FULL_THRESHOLD(7)
      )
     pcie_4_0_512b_async_fifo_blk
       (
    // Write side
    .clk_i(user_clk2_i),
    .clk_en_i(user_clk_en_i),
        .reset_n_i(reset_n_user_clk2_i),
        .link_down_reset_i(link_down_reset_i),
    .write_data_i(fifo_in_data),
    .write_en_i(fifo_in_data_valid),
    .fifo_almost_full_o(fifo_almost_full_user_clk),
    // Read side
    .read_en_i(output_mux_ready),
    .read_data_o(fifo_read_data),
    .read_data_valid_o(fifo_read_data_valid)
    );

   // Instance of output MUX
   xp4_usp_smsw_512b_cc_output_mux #
     (
      .TCQ(TCQ),
      .IMPL_TARGET(IMPL_TARGET),
      .IN_DATA_WIDTH(OUTPUT_MUX_IN_DATA_WIDTH),
      .OUT_DATA_WIDTH(AXI4_CORE_DATA_WIDTH),
      .TUSER_WIDTH(AXI4_CORE_CC_TUSER_WIDTH),
      .TKEEP_WIDTH(AXI4_CORE_CC_TKEEP_WIDTH),
      .TREADY_WIDTH(AXI4_CORE_CC_TREADY_WIDTH)
      )
     pcie_4_0_512b_cc_output_mux_blk
       (
        .clk_i(user_clk2_i),
        .reset_n_i(reset_n_user_clk2_i),
        .link_down_reset_i(link_down_reset_i),
    .in_data_i(fifo_read_data),
    .in_data_valid_i(fifo_read_data_valid),
    .upstream_ready_o(output_mux_ready),

    .out_data_o(core_cc_tdata_o),
        .out_data_valid_o(core_cc_tvalid_o),
    .out_tuser_o(core_cc_tuser_o),
    .out_tlast_o(core_cc_tlast_o),
    .out_tkeep_o(core_cc_tkeep_o),
    .downstream_ready_i(core_cc_tready_int)
    );


endmodule // pcie4_0_512b_cc_intfc







   
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_512b_cc_output_mux.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_512b_cc_output_mux #(
   parameter TCQ = 100,
   parameter IMPL_TARGET = "SOFT",
   parameter IN_DATA_WIDTH = 256+33+8+1,    
   parameter OUT_DATA_WIDTH = 256,
   parameter TUSER_WIDTH = 33,
   parameter TKEEP_WIDTH = 8,
   parameter TREADY_WIDTH = 4
   )
  (
    input  wire           clk_i // 500 MHz clock for core-facing interfaces
   ,input  wire           reset_n_i // Reset in the user clock domain
   ,input  wire           link_down_reset_i // Link went down

   ,input wire[IN_DATA_WIDTH-1:0] in_data_i
   ,input wire in_data_valid_i
   ,output wire upstream_ready_o

   ,output reg [OUT_DATA_WIDTH-1:0]  out_data_o
   ,output reg           out_data_valid_o
   ,output reg [TUSER_WIDTH-1:0] out_tuser_o
   ,output reg          out_tlast_o
   ,output reg [TKEEP_WIDTH-1:0] out_tkeep_o
   ,input  wire [TREADY_WIDTH-1:0]  downstream_ready_i
   );


   reg [1:0] output_fifo_occupancy;
  reg          output_fifo_write_ptr;
  reg          output_fifo_read_ptr;
   wire      output_fifo_full;
   wire      output_fifo_empty;

   reg [OUT_DATA_WIDTH-1:0] m_axis_cc_tdata_first_reg;
   reg [TKEEP_WIDTH-1:0]    m_axis_cc_tkeep_first_reg;
   reg [TUSER_WIDTH-1:0]    m_axis_cc_tuser_first_reg;
   reg                 m_axis_cc_tlast_first_reg;
   
   reg [OUT_DATA_WIDTH-1:0] m_axis_cc_tdata_second_reg;
   reg [TKEEP_WIDTH-1:0]    m_axis_cc_tkeep_second_reg;
   reg [TUSER_WIDTH-1:0]    m_axis_cc_tuser_second_reg;
   reg                 m_axis_cc_tlast_second_reg;
   
   wire             output_reg_mux_sel;
   //---------------------------------------------------------------------------------------------
   // Output FIFO.
   // The main FIFO feeds into two read registers in the core clock domain, which are configured
   // as a 2-entry FIFO.
   // This can be thought of as logical extensions of the main FIFO.
   //---------------------------------------------------------------------------------------------

   assign    upstream_ready_o = ~output_fifo_full;

   // Maintain write and read pointers
   always @(posedge clk_i)
     if (~reset_n_i)
       output_fifo_write_ptr <= #(TCQ)  1'b0;
     else if (link_down_reset_i)
       output_fifo_write_ptr <= #(TCQ)  1'b0;
     else
       if (in_data_valid_i & ~output_fifo_full)
     output_fifo_write_ptr <= #(TCQ) ~output_fifo_write_ptr;
   
   always @(posedge clk_i)
     if (~reset_n_i)
       output_fifo_read_ptr <= #(TCQ) 2'd0;
     else if (link_down_reset_i)
       output_fifo_read_ptr <= #(TCQ) 2'd0;
     else
       if ((downstream_ready_i[3] | ~out_data_valid_o) &
       ~output_fifo_empty)
     output_fifo_read_ptr <= #(TCQ) ~output_fifo_read_ptr;

      // Maintain FIFO occupancy
   always @(posedge clk_i)
     if (~reset_n_i)
       output_fifo_occupancy <= #(TCQ)  2'd0;
     else if (link_down_reset_i)
       output_fifo_occupancy <= #(TCQ)  2'd0;
     else
       if ((in_data_valid_i & ~output_fifo_full) &
       ~((downstream_ready_i[3] | ~out_data_valid_o) &
         ~output_fifo_empty))
     output_fifo_occupancy <= #(TCQ) output_fifo_occupancy + 2'd1;
       else
     if (~(in_data_valid_i & ~output_fifo_full) &
         ((downstream_ready_i[3] | ~out_data_valid_o) &
          ~output_fifo_empty))
       output_fifo_occupancy <= #(TCQ) output_fifo_occupancy - 2'd1;
   
   assign output_fifo_full = output_fifo_occupancy[1];
   assign output_fifo_empty = (output_fifo_occupancy == 2'b00);

   // Write data into the Output registers
   always @(posedge clk_i)
     if (~reset_n_i)
       begin
          m_axis_cc_tdata_first_reg <= #(TCQ) {OUT_DATA_WIDTH{1'b0}};
          m_axis_cc_tdata_second_reg <= #(TCQ) {OUT_DATA_WIDTH{1'b0}};
          m_axis_cc_tkeep_first_reg <= #(TCQ) {TKEEP_WIDTH{1'b0}};
          m_axis_cc_tkeep_second_reg <= #(TCQ) {TKEEP_WIDTH{1'b0}};
          m_axis_cc_tuser_first_reg <= #(TCQ) {TUSER_WIDTH{1'b0}};
          m_axis_cc_tuser_second_reg <= #(TCQ) {TUSER_WIDTH{1'b0}};
          m_axis_cc_tlast_first_reg <= #(TCQ) 1'b0;
          m_axis_cc_tlast_second_reg <= #(TCQ) 1'b0;
       end
     else
        if (in_data_valid_i & ~output_fifo_full)
      begin
        case(output_fifo_write_ptr)
          1'b0:
         begin
            m_axis_cc_tdata_first_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH-1:0];
            m_axis_cc_tkeep_first_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH-1:OUT_DATA_WIDTH];
            m_axis_cc_tuser_first_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH+TUSER_WIDTH-1:OUT_DATA_WIDTH+TKEEP_WIDTH];
            m_axis_cc_tlast_first_reg <= #(TCQ) in_data_i[IN_DATA_WIDTH-1];
         end
           default:
         begin
            m_axis_cc_tdata_second_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH-1:0];
            m_axis_cc_tkeep_second_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH-1:OUT_DATA_WIDTH];
            m_axis_cc_tuser_second_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH+TUSER_WIDTH-1:OUT_DATA_WIDTH+TKEEP_WIDTH];
            m_axis_cc_tlast_second_reg <= #(TCQ) in_data_i[IN_DATA_WIDTH-1];
         end
         endcase // case(output_fifo_write_ptr)
        end // if (in_data_valid_i & ~output_fifo_full)
   
   // Output registers

   assign output_reg_mux_sel = output_fifo_read_ptr;

   always @(posedge clk_i)
     if (~reset_n_i)
       begin
      out_data_o <= #(TCQ)  {OUT_DATA_WIDTH{1'b0}};
      out_tuser_o <= #(TCQ)  {TUSER_WIDTH{1'b0}};
      out_tkeep_o <= #(TCQ)  {TKEEP_WIDTH{1'b0}};
      out_tlast_o <= #(TCQ)  1'b0;
       end
     else
       begin
      if (~out_data_valid_o | downstream_ready_i[0])
        begin
           case(output_reg_mux_sel)
         1'b0:
           begin
              out_data_o[127:0] <= #(TCQ)  m_axis_cc_tdata_first_reg[127:0];
           end
         default:
           begin
              out_data_o[127:0] <= #(TCQ)  m_axis_cc_tdata_second_reg[127:0];
           end
           endcase // case(output_reg_mux_sel)
        end // if (~out_data_valid_o | downstream_ready_i[0])

      if (~out_data_valid_o | downstream_ready_i[1])
        begin
           case(output_reg_mux_sel)
         1'b0:
           begin
              out_data_o[255:128] <= #(TCQ)  m_axis_cc_tdata_first_reg[255:128];
           end
         default:
           begin
              out_data_o[255:128] <= #(TCQ)  m_axis_cc_tdata_second_reg[255:128];
           end
           endcase // case(output_reg_mux_sel)
        end // if (~out_data_valid_o | downstream_ready_i[1])
      
      if (~out_data_valid_o | downstream_ready_i[2])
        begin
           case(output_reg_mux_sel)
         1'b0:
           begin
              out_tuser_o <= #(TCQ)  m_axis_cc_tuser_first_reg;
           end
         default:
           begin
              out_tuser_o <= #(TCQ)  m_axis_cc_tuser_second_reg;
           end
           endcase // case(output_reg_mux_sel)
        end // if (~out_data_valid_o | downstream_ready_i[2])
      
      if (~out_data_valid_o | downstream_ready_i[3])
        begin
           case(output_reg_mux_sel)
         1'b0:         
           begin
              out_tkeep_o <= #(TCQ)  m_axis_cc_tkeep_first_reg;
              out_tlast_o <= #(TCQ)  m_axis_cc_tlast_first_reg;
           end
         default:
           begin
              out_tkeep_o <= #(TCQ)  m_axis_cc_tkeep_second_reg;
              out_tlast_o <= #(TCQ)  m_axis_cc_tlast_second_reg;
           end
           endcase // case(output_reg_mux_sel)
        end // if (~out_data_valid_o | downstream_ready_i[3])
       end // else: !if(~reset_n_i)

   always @(posedge clk_i)
     if (~reset_n_i)
       out_data_valid_o <= #(TCQ) 1'b0;
     else
       if (~out_data_valid_o | downstream_ready_i[0])
     out_data_valid_o <= #(TCQ) ~output_fifo_empty;

endmodule // pcie_4_0_512b_cc_output_mux

//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_512b_cq_intfc.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_512b_cq_intfc #(
   parameter TCQ = 100,
   parameter IMPL_TARGET = "SOFT",
   parameter AXISTEN_IF_EXT_512_INTFC_RAM_STYLE = "SRL",
   parameter AXI4_USER_DATA_WIDTH = 512,
   parameter AXI4_CORE_DATA_WIDTH = 256,
   parameter AXI4_USER_CQ_TUSER_WIDTH = 183,
   parameter AXI4_CORE_CQ_TUSER_WIDTH = 88,
   parameter AXI4_USER_CQ_TKEEP_WIDTH = 16,
   parameter AXI4_CORE_CQ_TKEEP_WIDTH = 8,
   parameter AXI4_CORE_CQ_TREADY_WIDTH = 22,
   parameter PARITY_ENABLE = 0
   ) 
  (
    input  wire           user_clk2_i // 500 MHz clock for core-facing interfaces
   ,input  wire           user_clk_i // 250 MHz clock for client-facing interfaces
   ,input  wire           user_clk_en_i // User clock enable for clock domain crossing
   ,input  wire           reset_n_user_clk_i // Reset in the user clock domain
   ,input  wire           reset_n_user_clk2_i // Reset in the user clock2 domain
   ,input  wire           link_down_reset_i // Link went down
   // Attributes
   ,input  wire           attr_straddle_en_i // Enable straddle
   ,input wire [1:0]      attr_alignment_mode_i // Payload alignment mode
                                                // (00= Dword-aligned, 10 = 128b address-aligned)
   //-----------------------------------------------------------------------------------------------
   // Client-side signals
   //-----------------------------------------------------------------------------------------------
   ,output wire [AXI4_USER_DATA_WIDTH-1:0]   m_axis_cq_tdata_o
   ,output wire           m_axis_cq_tvalid_o
   ,output wire [AXI4_USER_CQ_TUSER_WIDTH-1:0]   m_axis_cq_tuser_o
   ,output wire           m_axis_cq_tlast_o
   ,output wire [AXI4_USER_CQ_TKEEP_WIDTH-1:0]    m_axis_cq_tkeep_o
   ,input  wire           m_axis_cq_tready_i
   ,input  wire [1:0]     pcie_cq_np_req_i // Client request to deliver NP TLP
   ,output wire [5:0]     pcie_cq_np_req_count_o // Current value of interface credit count for NP TLPs
   //-----------------------------------------------------------------------------------------------
   // Core-side signals
   //-----------------------------------------------------------------------------------------------
   ,input  wire [AXI4_CORE_DATA_WIDTH-1:0] core_cq_tdata_i
   ,input  wire           core_cq_tvalid_i
   ,input  wire [AXI4_CORE_CQ_TUSER_WIDTH-1:0] core_cq_tuser_i
   ,input  wire           core_cq_tlast_i
   ,input  wire [AXI4_CORE_CQ_TKEEP_WIDTH-1:0] core_cq_tkeep_i
   ,output wire [AXI4_CORE_CQ_TREADY_WIDTH-1:0] core_cq_tready_o
   ,output reg            posted_req_delivered_o // Signals the delivery of a Posted Req on the CQ interface
   ,output reg            cq_pipeline_empty_o // Indicates that the entire CQ pipeline of the bridge is empty.
   ,output reg            cq_np_user_credit_rcvd_o // Indicates that the user issued one NP credit
   );

   localparam FIFO_WIDTH = PARITY_ENABLE? (AXI4_CORE_DATA_WIDTH + AXI4_CORE_CQ_TUSER_WIDTH + 
                       AXI4_CORE_CQ_TKEEP_WIDTH + 1)*2 +2 :
               (AXI4_CORE_DATA_WIDTH + AXI4_CORE_CQ_TUSER_WIDTH + 
                AXI4_CORE_CQ_TKEEP_WIDTH + 1)*2 +2 -64;

   localparam TUSER_LOWER_OFFSET = AXI4_CORE_DATA_WIDTH + AXI4_CORE_CQ_TKEEP_WIDTH;
   localparam TUSER_UPPER_OFFSET = PARITY_ENABLE? AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_CQ_TKEEP_WIDTH*2 +
                   AXI4_CORE_CQ_TUSER_WIDTH +2:
                   AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_CQ_TKEEP_WIDTH*2 +
                   AXI4_CORE_CQ_TUSER_WIDTH +2 -32;
   
  localparam FIFO_READ_DATA_UPPER_OFFSET = PARITY_ENABLE?
                   AXI4_CORE_DATA_WIDTH + AXI4_CORE_CQ_TKEEP_WIDTH + AXI4_CORE_CQ_TUSER_WIDTH +2:
                   AXI4_CORE_DATA_WIDTH + AXI4_CORE_CQ_TKEEP_WIDTH + AXI4_CORE_CQ_TUSER_WIDTH +2 -32;
  
  localparam FIFO_READ_TKEEP_UPPER_OFFSET = PARITY_ENABLE?
                    AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_CQ_TKEEP_WIDTH + AXI4_CORE_CQ_TUSER_WIDTH +2:
                                    AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_CQ_TKEEP_WIDTH + AXI4_CORE_CQ_TUSER_WIDTH +2 -32;

   localparam OUTPUT_MUX_IN_DATA_WIDTH = AXI4_USER_DATA_WIDTH +
                     AXI4_USER_CQ_TKEEP_WIDTH +
                     AXI4_USER_CQ_TUSER_WIDTH + 1;

   (* KEEP = "true" *) reg [AXI4_CORE_CQ_TREADY_WIDTH-1:0] core_cq_tready_reg;
   (* KEEP = "true" *) reg core_cq_tready_user_clk2;

   reg [AXI4_CORE_DATA_WIDTH-1:0] core_cq_tdata_reg_upper;
   reg [AXI4_CORE_DATA_WIDTH-1:0] core_cq_tdata_reg_lower;
   reg [AXI4_CORE_CQ_TUSER_WIDTH-1:0] core_cq_tuser_reg_upper;
   reg [AXI4_CORE_CQ_TUSER_WIDTH-1:0] core_cq_tuser_reg_lower;
   reg                       core_cq_tlast_reg_upper;
   reg                       core_cq_tlast_reg_lower;
   reg [AXI4_CORE_CQ_TKEEP_WIDTH-1:0] core_cq_tkeep_reg_upper;
   reg [AXI4_CORE_CQ_TKEEP_WIDTH-1:0] core_cq_tkeep_reg_lower;
   reg                       core_cq_tvalid_reg_upper;
   reg                       core_cq_tvalid_reg_lower;

   wire                   fifo_almost_full_user_clk;

   wire [FIFO_WIDTH-1:0]           fifo_in_data;
   reg [FIFO_WIDTH-1:0]           fifo_in_data_reg;
   reg                       fifo_in_data_valid_reg;
   reg                       fifo_read_en;
   wire                   fifo_read_data_valid;
   wire [FIFO_WIDTH-1:0]           fifo_read_data;

   wire [3:0]                   read_first_be_lower;
   wire [3:0]                   read_last_be_lower;
   wire [31:0]                   read_byte_en_lower;
   wire                   read_sop_lower;
   wire                   read_discontinue_lower;
   wire                   read_tph_present_lower;
   wire [1:0]                   read_tph_type_lower;
   wire [7:0]                   read_tph_st_tag_lower;
   wire [2:0]                   read_eop_ptr_lower;
   wire                   read_tlast_lower;
   wire                   read_tlast_upper;
   wire                   read_data_valid_lower;
   wire                   read_data_valid_upper;

   wire [3:0]                   read_first_be_upper;
   wire [3:0]                   read_last_be_upper;
   wire [31:0]                   read_byte_en_upper;
   wire                   read_sop_upper;
   wire                   read_discontinue_upper;
   wire                   read_tph_present_upper;
   wire [1:0]                   read_tph_type_upper;
   wire [7:0]                   read_tph_st_tag_upper;
   wire [2:0]                   read_eop_ptr_upper;

   reg [1:0]                   read_data_valid_reg;
   reg [FIFO_WIDTH-1:0]           read_data_reg;
   reg [FIFO_WIDTH/2-1:0]           saved_data_reg;
   reg                       saved_eop;
   reg                       saved_err;
   
   wire [3:0]                   read_data_reg_first_be_lower;
   wire [3:0]                   read_data_reg_last_be_lower;
   wire [31:0]                   read_data_reg_byte_en_lower;
   wire                    read_data_reg_sop_lower;
   wire                    read_data_reg_discontinue_lower;
   wire                    read_data_reg_tph_present_lower;
   wire [1:0]                   read_data_reg_tph_type_lower;
   wire [7:0]                   read_data_reg_tph_st_tag_lower;
   wire [31:0]                   read_data_reg_parity_lower;
   wire [2:0]                   read_data_reg_eop_ptr_lower;
   wire [3:0]                   read_data_reg_first_be_upper;
   wire [3:0]                   read_data_reg_last_be_upper;
   wire [31:0]                   read_data_reg_byte_en_upper;
   wire                    read_data_reg_sop_upper;
   wire                    read_data_reg_discontinue_upper;
   wire                    read_data_reg_tph_present_upper;
   wire [1:0]                   read_data_reg_tph_type_upper;
   wire [7:0]                   read_data_reg_tph_st_tag_upper;
   wire [31:0]                   read_data_reg_parity_upper;
   wire [2:0]                   read_data_reg_eop_ptr_upper;
  wire                       read_data_reg_tlast_lower;
  wire                       read_data_reg_tlast_upper;
   wire                   sop_in_lower_half;
   wire                   sop_in_upper_half;
   wire                   eop_in_lower_half;
   wire                   eop_in_upper_half;

   wire [7:0]                   read_data_out_first_be;
   wire [7:0]                   read_data_out_last_be;
   wire [63:0]                   read_data_out_byte_en;
   wire [1:0]                   read_data_out_is_sop;
   wire [1:0]                   read_data_out_is_sop0_ptr;
   wire [1:0]                   read_data_out_is_sop1_ptr;
   wire [1:0]                   read_data_out_is_eop;
   wire [3:0]                   read_data_out_is_eop0_ptr;
   wire [3:0]                   read_data_out_is_eop1_ptr;
   wire                   read_data_out_discontinue;
   wire [1:0]                   read_data_out_tph_present;
   wire [3:0]                   read_data_out_tph_type;
   wire [15:0]                   read_data_out_tph_st_tag;
   wire [63:0]                   read_data_out_parity;
   
   wire [ AXI4_USER_CQ_TUSER_WIDTH-1:0] read_data_out_tuser;
   wire [ AXI4_USER_DATA_WIDTH-1:0]     read_data_out_tdata;
   wire [ AXI4_USER_CQ_TKEEP_WIDTH-1:0] read_data_out_tkeep;
   wire                 read_data_out_tlast;
   
   wire [OUTPUT_MUX_IN_DATA_WIDTH-1:0]     output_mux_in_data;

   wire                 output_mux_ready;
   
   wire [1:0]                 cq_np_user_credit_rcvd_user_clk;
   wire [1:0]                 posted_req_delivered_user_clk;

   wire                 pipeline_empty_user_clk;
   wire                 out_mux_pipeline_empty;
   reg                     pipeline_empty_core_clk;
   reg [2:0]                 cq_pipeline_empty_reg;

   // Read State Machine states
   localparam                           IDLE = 2'd0;
   localparam                           EXPECT_NEW_WORD = 2'd1;
   localparam                           SEND_SAVED_HALF_WORD = 2'd2;
   localparam                           WAIT_FOR_UPPER_HALF = 2'd3;
   reg [1:0]                 read_state;

   // Capture incoming data from core at 500 MHz into upper and lower registers
   always @(posedge user_clk2_i)
     if (~reset_n_user_clk2_i)
       begin
      core_cq_tdata_reg_upper <= #TCQ {AXI4_CORE_DATA_WIDTH{1'b0}};
      core_cq_tdata_reg_lower <= #TCQ {AXI4_CORE_DATA_WIDTH{1'b0}};
      core_cq_tuser_reg_upper <= #TCQ {AXI4_CORE_CQ_TUSER_WIDTH{1'b0}};
      core_cq_tuser_reg_lower <= #TCQ {AXI4_CORE_CQ_TUSER_WIDTH{1'b0}};
      core_cq_tkeep_reg_upper <= #TCQ {AXI4_CORE_CQ_TKEEP_WIDTH{1'b0}};
      core_cq_tkeep_reg_lower <= #TCQ {AXI4_CORE_CQ_TKEEP_WIDTH{1'b0}};
      core_cq_tlast_reg_upper <= #TCQ 1'b0;
      core_cq_tlast_reg_lower <= #TCQ 1'b0;
       core_cq_tvalid_reg_upper <= #TCQ 1'b0;
      core_cq_tvalid_reg_lower <= #TCQ 1'b0;
       end // if (~reset_n_user_clk_i)
     else
       if (user_clk_en_i)
     begin
        core_cq_tdata_reg_lower <= #TCQ core_cq_tdata_i;
        core_cq_tuser_reg_lower <= #TCQ core_cq_tuser_i;
        core_cq_tkeep_reg_lower <= #TCQ core_cq_tkeep_i;
        core_cq_tlast_reg_lower <= #TCQ core_cq_tlast_i;
        core_cq_tvalid_reg_lower <= #TCQ core_cq_tvalid_i & core_cq_tready_user_clk2;
     end
       else
     begin
        core_cq_tdata_reg_upper <= #TCQ core_cq_tdata_i;
        core_cq_tuser_reg_upper <= #TCQ core_cq_tuser_i;
        core_cq_tkeep_reg_upper <= #TCQ core_cq_tkeep_i;
        core_cq_tlast_reg_upper <= #TCQ core_cq_tlast_i;
        core_cq_tvalid_reg_upper <= #TCQ core_cq_tvalid_i & core_cq_tready_user_clk2;
     end // else: !if(user_clk_en_i)

   // Write data into FIFO using 250 MHz user_clk

  generate
    if (PARITY_ENABLE)
      assign fifo_in_data =
          {
       core_cq_tvalid_reg_upper,
       core_cq_tlast_reg_upper,
       core_cq_tuser_reg_upper,
       core_cq_tkeep_reg_upper,
       core_cq_tdata_reg_upper,
       core_cq_tvalid_reg_lower,
       core_cq_tlast_reg_lower,
       core_cq_tuser_reg_lower,
       core_cq_tkeep_reg_lower,
       core_cq_tdata_reg_lower
       };
    else
      assign fifo_in_data =
          {
       core_cq_tvalid_reg_upper,
       core_cq_tlast_reg_upper,
       core_cq_tuser_reg_upper[87:85],
       core_cq_tuser_reg_upper[52:0],
       core_cq_tkeep_reg_upper,
       core_cq_tdata_reg_upper,
       core_cq_tvalid_reg_lower,
       core_cq_tlast_reg_lower,
       core_cq_tuser_reg_lower[87:85],
       core_cq_tuser_reg_lower[52:0],
       core_cq_tkeep_reg_lower,
       core_cq_tdata_reg_lower
       };
  endgenerate

   always @(posedge user_clk_i)
     if (~reset_n_user_clk_i)
       begin
      fifo_in_data_reg <= #TCQ {FIFO_WIDTH{1'b0}};      
      fifo_in_data_valid_reg <= #TCQ 1'b0;
       end
     else
       begin
      fifo_in_data_reg <= #TCQ fifo_in_data;
         fifo_in_data_valid_reg <= #TCQ (core_cq_tvalid_reg_lower |
                     core_cq_tvalid_reg_upper);
       end // else: !if(~reset_n_user_clk_i)

   // Generate ready to core in the user_clk2 domain
   always @(posedge user_clk2_i)
     if (~reset_n_user_clk2_i)
       begin
      core_cq_tready_user_clk2 <= #TCQ 1'b0;
      core_cq_tready_reg <= #TCQ {AXI4_CORE_CQ_TREADY_WIDTH{1'b0}};
       end
     else
       begin
             core_cq_tready_user_clk2 <= #TCQ ~fifo_almost_full_user_clk;
      core_cq_tready_reg <= #TCQ {AXI4_CORE_CQ_TREADY_WIDTH{~fifo_almost_full_user_clk}};
       end

   assign core_cq_tready_o = core_cq_tready_reg;
   
   // Main FIFO instance
   xp4_usp_smsw_512b_sync_fifo #
     (
      .TCQ(TCQ),
      .IMPL_TARGET(IMPL_TARGET),
      .AXISTEN_IF_EXT_512_INTFC_RAM_STYLE(AXISTEN_IF_EXT_512_INTFC_RAM_STYLE),
      .FIFO_WIDTH(FIFO_WIDTH),
      .FIFO_DEPTH(8),
      .FIFO_ALMOST_FULL_THRESHOLD(5)
      )
     pcie_4_0_512b_sync_fifo_blk
       (
        .clk_i(user_clk_i),
        .reset_n_i(reset_n_user_clk_i),
        .link_down_reset_i(link_down_reset_i),
    .write_data_i(fifo_in_data_reg),
    .write_en_i(fifo_in_data_valid_reg),
    .read_en_i(fifo_read_en),
    .read_data_o(fifo_read_data),
    .read_data_valid_o(fifo_read_data_valid),
    .fifo_almost_full(fifo_almost_full_user_clk)
    );
   
   // Read-side logic
   
   assign read_first_be_lower = fifo_read_data[TUSER_LOWER_OFFSET +3:
                           TUSER_LOWER_OFFSET];
   assign read_last_be_lower = fifo_read_data[TUSER_LOWER_OFFSET +7:
                          TUSER_LOWER_OFFSET +4];
   assign read_byte_en_lower = fifo_read_data[TUSER_LOWER_OFFSET +39:
                             TUSER_LOWER_OFFSET +8];
   assign read_sop_lower = fifo_read_data[TUSER_LOWER_OFFSET + 40];
   assign read_discontinue_lower = fifo_read_data[TUSER_LOWER_OFFSET + 41];
   assign read_tph_present_lower = fifo_read_data[TUSER_LOWER_OFFSET + 42];  
   assign read_tph_type_lower = fifo_read_data[TUSER_LOWER_OFFSET + 44:
                        TUSER_LOWER_OFFSET + 43];
   assign read_tph_st_tag_lower = fifo_read_data[TUSER_LOWER_OFFSET + 52:   
                            TUSER_LOWER_OFFSET + 45];
  generate
    if (PARITY_ENABLE)
      assign read_eop_ptr_lower = fifo_read_data[TUSER_LOWER_OFFSET + 87:
                         TUSER_LOWER_OFFSET + 85];
    else
      assign read_eop_ptr_lower = fifo_read_data[TUSER_LOWER_OFFSET + 55:
                         TUSER_LOWER_OFFSET + 53];
  endgenerate


  assign     read_first_be_upper = fifo_read_data[TUSER_UPPER_OFFSET +3:
                           TUSER_UPPER_OFFSET];
   assign read_last_be_upper = fifo_read_data[TUSER_UPPER_OFFSET +7:
                          TUSER_UPPER_OFFSET +4];
   assign read_byte_en_upper = fifo_read_data[TUSER_UPPER_OFFSET +39:
                             TUSER_UPPER_OFFSET +8];
   assign read_sop_upper = fifo_read_data[TUSER_UPPER_OFFSET + 40];
   assign read_discontinue_upper = fifo_read_data[TUSER_UPPER_OFFSET + 41];
   assign read_tph_present_upper = fifo_read_data[TUSER_UPPER_OFFSET + 42];  
   assign read_tph_type_upper = fifo_read_data[TUSER_UPPER_OFFSET + 44:
                        TUSER_UPPER_OFFSET + 43];
   assign read_tph_st_tag_upper = fifo_read_data[TUSER_UPPER_OFFSET + 52:   
                            TUSER_UPPER_OFFSET + 45];
  generate
    if (PARITY_ENABLE)
      assign read_eop_ptr_upper = fifo_read_data[TUSER_UPPER_OFFSET + 87:
                         TUSER_UPPER_OFFSET + 85];
    else
      assign read_eop_ptr_upper = fifo_read_data[TUSER_UPPER_OFFSET + 55:
                           TUSER_UPPER_OFFSET + 53];
  endgenerate

  generate
    if (PARITY_ENABLE)
      begin
    assign     read_tlast_lower = fifo_read_data[AXI4_CORE_DATA_WIDTH + AXI4_CORE_CQ_TKEEP_WIDTH +
                             AXI4_CORE_CQ_TUSER_WIDTH];
    assign     read_tlast_upper = fifo_read_data[AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_CQ_TKEEP_WIDTH*2 +
                             AXI4_CORE_CQ_TUSER_WIDTH*2 +2];
      end
    else
      begin
    assign     read_tlast_lower = fifo_read_data[AXI4_CORE_DATA_WIDTH + AXI4_CORE_CQ_TKEEP_WIDTH +
                             AXI4_CORE_CQ_TUSER_WIDTH -32];
    assign     read_tlast_upper = fifo_read_data[AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_CQ_TKEEP_WIDTH*2 +
                             AXI4_CORE_CQ_TUSER_WIDTH*2 +2 -64];
      end // else: !if(PARITY_ENABLE)
  endgenerate

    assign        read_data_valid_lower = fifo_read_data[FIFO_WIDTH/2-1] & fifo_read_data_valid;
    assign        read_data_valid_upper = fifo_read_data[FIFO_WIDTH-1] & fifo_read_data_valid;


   // Read State Machine States
   //
   // IDLE: Currently not forwarding a packet.  Read data register is either empty, or contains the last beat of a packet.
   // EXPECT_NEW_WORD: Currently forwarding a packet, and there is no data saved from a previous beat
   // SEND_SAVED_HALF_WORD: There is a half-word saved from a previous beat in the saved data register.
   // WAIT_FOR_UPPER_HALF: There is a half-word saved from a previous beat in the read data register which does not end with an EOP.
   
   always @(posedge user_clk_i)
     if (~reset_n_user_clk_i)
       begin
      read_data_valid_reg <= #TCQ 2'b00;
      read_state <= #TCQ IDLE;
       end
     else if (link_down_reset_i)
       begin
      read_data_valid_reg <= #TCQ 2'b00;
      read_state <= #TCQ IDLE;
       end
     else
    case(read_state)
      IDLE:
        begin
           // IDLE: Currently not forwarding a packet.  Read data register is either empty, or contains the last beat of a packet.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if (read_data_valid_lower)
              // New TLP starting in the lower half of the incoming word.
              // Update the lower half of the data register with the lower half of the incoming word.
              begin
             if (read_data_valid_upper)
               // Both halves of the incoming word have valid data in them.
               begin
                  // If straddle is not enabled and the packet in the upper half is a new one,
                  // Save it for next cycle.
                  // Also, if the packet in the lower half ends with an error, do not fill the upper half.
                  if ((~attr_straddle_en_i & read_sop_upper)|
                  read_discontinue_lower)
                begin
                   read_data_valid_reg <= #TCQ 2'b01;
                   read_state <= #TCQ SEND_SAVED_HALF_WORD;
                end
                  else
                begin
                   read_data_valid_reg <= #TCQ 2'b11;
                   if (read_tlast_upper)
                     read_state <= #TCQ IDLE;
                   else
                     read_state <= #TCQ EXPECT_NEW_WORD;
                end // else: !if(~attr_straddle_en_i & read_sop_upper)
               end // if (read_data_valid_upper)
             else
               begin
                  // New TLP started in the lower half, but there is no valid data in the upper half.
                  if (read_tlast_lower)
                // We have a complete TLP in the lower half, send it.
                begin
                   read_data_valid_reg <= #TCQ 2'b01;
                   read_state <= #TCQ IDLE;
                end
                  else
                begin
                   // Wait for more data to fill upper half of read data register.
                   read_data_valid_reg <= #TCQ 2'b00;
                   read_state <= #TCQ WAIT_FOR_UPPER_HALF;
                end // else: !if(read_tlast_lower)
               end // else: !if(read_data_valid_upper)
              end // if (read_data_valid_lower)
            else
              if (read_data_valid_upper)
            begin
               // No valid data in the lower half of the incoming word, but there is a packet starting in the upper half.
               if (read_tlast_upper)
                 // We have a complete packet, send it in the lower half.
                 begin
                read_data_valid_reg <= #TCQ 2'b01;
                read_state <= #TCQ IDLE;
                 end
               else
                 begin
                // Save the upper half of the incoming word
                // and wait for more data.
                read_data_valid_reg <= #TCQ 2'b00;
                read_state <= #TCQ WAIT_FOR_UPPER_HALF;
                 end // else: !if(read_tlast_upper)
            end // if (read_data_valid_upper)
              else
            // No valid data from FIFO
            begin
               if (output_mux_ready)
                 read_data_valid_reg <= #TCQ 2'b00;
               read_state <= #TCQ IDLE;
            end // else: !if(read_data_valid_upper)
         end // if ((read_data_valid_reg == 2'b00) | output_mux_ready)
        end // case: IDLE
      
      EXPECT_NEW_WORD:
        begin
           // Currently forwarding a packet.  There is no saved data.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if (read_data_valid_lower)
              // New data starting in the lower half of the incoming word.
              // Update the lower half of the data register with the lower half of the incoming word.
              begin
             if (read_data_valid_upper)
               // Both halves of the incoming word have valid data in them.
               begin
                  // If straddle is not enabled and the packet in the upper half is a new one,
                  // Save it for next cycle.
                  // Also, if the packet in the lower half ends with an error, do not fill the upper half.
                  if ((~attr_straddle_en_i & read_sop_upper)|
                  read_discontinue_lower)
                begin
                   read_data_valid_reg <= #TCQ 2'b01;
                   read_state <= #TCQ SEND_SAVED_HALF_WORD;
                end
                  else
                begin
                   read_data_valid_reg <= #TCQ 2'b11;
                   if (read_tlast_upper)
                     read_state <= #TCQ IDLE;
                   else
                     read_state <= #TCQ EXPECT_NEW_WORD;
                end // else: !if(~attr_straddle_en_i & read_sop_upper)
               end // if (read_data_valid_upper)
             else
               begin
                  // Valid data in the lower half, but no valid data in the upper half.
                  if (read_tlast_lower)
                // We have the packet ending in the lower half, send it.
                begin
                   read_data_valid_reg <= #TCQ 2'b01;
                   read_state <= #TCQ IDLE;
                end
                  else
                begin
                   // Wait for more data to fill upper half of read data register.
                   read_data_valid_reg <= #TCQ 2'b00;
                   read_state <= #TCQ WAIT_FOR_UPPER_HALF;
                end // else: !if(read_tlast_lower)
               end // else: !if(read_data_valid_upper)
              end // if (read_data_valid_lower)
            else
              if (read_data_valid_upper)
            begin
               // No valid data in the lower half of the incoming word, but there is data in the upper half.
               if (read_tlast_upper)
                 // We have a complete packet, send it in the lower half.
                 begin
                read_data_valid_reg <= #TCQ 2'b01;
                read_state <= #TCQ IDLE;
                 end
               else
                 begin
                // Save the upper half of the incoming word
                // and wait for more data.
                read_data_valid_reg <= #TCQ 2'b00;
                read_state <= #TCQ WAIT_FOR_UPPER_HALF;
                 end // else: !if(read_tlast_upper)
            end // if (read_data_valid_upper)
              else
            // No valid data from FIFO
            begin
               if (output_mux_ready)
                 read_data_valid_reg <= #TCQ 2'b00;
               read_state <= #TCQ EXPECT_NEW_WORD;
            end // else: !if(read_data_valid_upper)
         end // if ((read_data_valid_reg == 2'b00) | output_mux_ready)
        end // case: EXPECT_NEW_WORD

      SEND_SAVED_HALF_WORD:
        begin
           // There is a half-word saved from a previous beat in the saved data register.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if ((~attr_straddle_en_i & saved_eop) | saved_err)
              // Saved data is the last beat of a packet and straddle is disabled.
              // Do not fill the upper half of read data register.
              begin
            read_data_valid_reg <= #TCQ 2'b01;
            read_state <= #TCQ IDLE;
              end
            else
              if (read_data_valid_lower)
            // New data starting in the lower half of the incoming word.
            // Update the upper half of the data register with the lower half of the incoming word.
            begin
               if (read_data_valid_upper)
                 // Both halves of the incoming word have valid data in them.
                 begin
                read_data_valid_reg <= #TCQ 2'b11;
                read_state <= #TCQ SEND_SAVED_HALF_WORD;
                 end
               else
                 begin
                read_data_valid_reg <= #TCQ 2'b11;
                if (read_tlast_lower)
                  read_state <= #TCQ IDLE;
                else
                  read_state <= #TCQ EXPECT_NEW_WORD;
                 end // else: !if(read_data_valid_upper)
            end // if (read_data_valid_lower)
              else
            if (read_data_valid_upper)
              begin
                 // No valid data in the lower half of the incoming word, but there is data in the upper half.
                 if (read_tlast_upper)
                   // We have a complete packet, send it in the upper half.
                   begin
                  read_data_valid_reg <= #TCQ 2'b11;
                  read_state <= #TCQ IDLE;
                   end
                 else
                   begin
                  read_data_valid_reg <= #TCQ 2'b11;
                  read_state <= #TCQ EXPECT_NEW_WORD;
                   end // else: !if(read_tlast_upper)
              end // if (read_data_valid_upper)
            else
              // No valid data from FIFO
              begin
                read_data_valid_reg <= #TCQ 2'b01;
                read_state <= #TCQ IDLE;
              end // else: !if(read_data_valid_upper)
         end // if ((read_data_valid_reg == 2'b00) | output_mux_ready)
        end // case: SEND_SAVED_HALF_WORD

      WAIT_FOR_UPPER_HALF:
        begin
           // There is a half-word saved from a previous beat in the read data register which does not end with an EOP.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if (read_data_valid_lower)
              // New data starting in the lower half of the incoming word.
              // Update the upper half of the data register with the lower half of the incoming word.
              begin
             read_data_valid_reg <= #TCQ 2'b11;
             if (read_data_valid_upper)
               // Both halves of the incoming word have valid data in them.
               begin
                 if (read_tlast_upper)
                   read_state <= #TCQ SEND_SAVED_HALF_WORD;
                 else
                   read_state <= #TCQ WAIT_FOR_UPPER_HALF;
               end
             else
               begin
                 if (read_tlast_lower)
                   read_state <= #TCQ IDLE;
                 else
                   read_state <= #TCQ EXPECT_NEW_WORD;
               end // else: !if(read_data_valid_upper)
              end // if (read_data_valid_lower)
            else
              if (read_data_valid_upper)
            begin
               // No valid data in the lower half of the incoming word, but there is data in the upper half.
               read_data_valid_reg <= #TCQ 2'b11;
               if (read_tlast_upper)
                 read_state <= #TCQ IDLE;
               else
                 read_state <= #TCQ EXPECT_NEW_WORD;
            end // if (read_data_valid_upper)
              else
            begin
               read_data_valid_reg <= #TCQ 2'b00;
               read_state <= #TCQ WAIT_FOR_UPPER_HALF;
            end // else: !if(read_data_valid_upper)
         end // if ((read_data_valid_reg == 2'b00) | output_mux_ready)
        end // case: WAIT_FOR_UPPER_HALF
    endcase // case(read_state)

   always @(posedge user_clk_i)
     if (~reset_n_user_clk_i)
       begin
      read_data_reg <= #TCQ {FIFO_WIDTH{1'b0}};
      saved_data_reg <= #TCQ {FIFO_WIDTH/2{1'b0}};
      saved_eop <= #TCQ 1'b0;
      saved_err <= #TCQ 1'b0;
       end
     else
    case(read_state)
      IDLE:
        begin
           // IDLE: Currently not forwarding a packet.  Read data register is either empty, or contains the last beat of a packet.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if (read_data_valid_lower)
              read_data_reg[FIFO_WIDTH/2-1:0] <= #TCQ fifo_read_data[FIFO_WIDTH/2-1:0];
            else
              read_data_reg[FIFO_WIDTH/2-1:0] <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
            read_data_reg[FIFO_WIDTH-1: FIFO_WIDTH/2] <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
            saved_data_reg <= #TCQ fifo_read_data[FIFO_WIDTH-1:FIFO_WIDTH/2];
            saved_eop <= #TCQ read_tlast_upper;
            saved_err <= #TCQ read_discontinue_upper;
         end
        end // case: IDLE

      EXPECT_NEW_WORD:
        begin
           // Currently not forwarding a packet.  
           // Read data register is either empty, or contains the last beat of a packet.           
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if (read_data_valid_lower)
              read_data_reg[FIFO_WIDTH/2-1:0] <= #TCQ fifo_read_data[FIFO_WIDTH/2-1:0];
            else
              read_data_reg[FIFO_WIDTH/2-1:0] <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
            read_data_reg[FIFO_WIDTH-1: FIFO_WIDTH/2] <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
            saved_data_reg <= #TCQ fifo_read_data[FIFO_WIDTH-1:FIFO_WIDTH/2];
            saved_eop <= #TCQ read_tlast_upper;
            saved_err <= #TCQ read_discontinue_upper;
         end
        end // case: EXPECT_NEW_WORD
      
      SEND_SAVED_HALF_WORD:
        begin
           // There is a half-word saved from a previous beat in the saved data register.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            read_data_reg[FIFO_WIDTH/2-1:0] <= #TCQ saved_data_reg[FIFO_WIDTH/2-1: 0];
            if (read_data_valid_lower)
              read_data_reg[FIFO_WIDTH-1: FIFO_WIDTH/2] <= #TCQ fifo_read_data[FIFO_WIDTH/2-1: 0];
            else
              read_data_reg[FIFO_WIDTH-1: FIFO_WIDTH/2] <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
            

            if ((~attr_straddle_en_i & saved_eop) | saved_err)
              // Save incoming data for next cycle.
              begin
             if (read_data_valid_lower)
               begin
                  saved_data_reg <= #TCQ fifo_read_data[FIFO_WIDTH/2-1: 0];
                  saved_eop <= #TCQ read_tlast_lower;
                  saved_err <= #TCQ read_discontinue_lower;
               end
             else
               begin
                  saved_data_reg <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
                  saved_eop <= #TCQ read_tlast_upper;
                  saved_err <= #TCQ read_discontinue_upper;
               end
              end
            else
              begin
             saved_data_reg <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
             saved_eop <= #TCQ read_tlast_upper;
             saved_err <= #TCQ read_discontinue_upper;
              end // else: !if((~attr_straddle_en_i & saved_eop) | saved_err)
         end // if ((read_data_valid_reg == 2'b00) | output_mux_ready)
        end // case: SEND_SAVED_HALF_WORD
      WAIT_FOR_UPPER_HALF:
        begin
           // There is a half-word saved from a previous beat in the read data register which does not end with an EOP.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
           read_data_reg[FIFO_WIDTH/2-1:0] <= #TCQ saved_data_reg[FIFO_WIDTH/2-1:0];
           if (read_data_valid_lower)
             read_data_reg[FIFO_WIDTH-1: FIFO_WIDTH/2] <= #TCQ fifo_read_data[FIFO_WIDTH/2-1: 0];
           else
             read_data_reg[FIFO_WIDTH-1: FIFO_WIDTH/2] <= #TCQ {FIFO_WIDTH/2{1'b0}};
             // Save incoming data for next cycle.
           saved_data_reg <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
           saved_eop <= #TCQ read_tlast_upper;
           saved_err <= #TCQ read_discontinue_upper;
         end
        end // case: WAIT_FOR_UPPER_HALF
    endcase // case(read_state)
         
   // Generate upstream ready
   always @(*)
     begin
    case(read_state)
      IDLE:
        begin
           fifo_read_en = (read_data_valid_reg == 2'b00) | output_mux_ready;
        end
      
      EXPECT_NEW_WORD:
        begin
           fifo_read_en = (read_data_valid_reg == 2'b00) | output_mux_ready;
        end

      SEND_SAVED_HALF_WORD:
        begin
           // There is a half-word saved from a previous beat in the saved data register.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if ((~attr_straddle_en_i & saved_eop) | saved_err)
              // Saved data is the last beat of a packet and straddle is disabled.
              // Do not fill the upper half of read data register.
              fifo_read_en = 1'b0;
            else
              fifo_read_en = 1'b1;
         end
           else
         fifo_read_en = 1'b0;
        end // case: SEND_SAVED_HALF_WORD

      WAIT_FOR_UPPER_HALF:
        begin
           // There is a half-word saved from a previous beat in the read data register which does not end with an EOP.
           fifo_read_en = (read_data_valid_reg == 2'b00) | output_mux_ready;
        end
    endcase // case(read_state)
     end // always @ (*)
   

   assign read_data_reg_first_be_lower = read_data_reg[TUSER_LOWER_OFFSET +3:
                               TUSER_LOWER_OFFSET];
   assign read_data_reg_last_be_lower = read_data_reg[TUSER_LOWER_OFFSET +7:
                              TUSER_LOWER_OFFSET +4];
   assign read_data_reg_byte_en_lower = read_data_reg[TUSER_LOWER_OFFSET +39:
                                 TUSER_LOWER_OFFSET +8];
   assign read_data_reg_sop_lower = read_data_reg[TUSER_LOWER_OFFSET + 40];
   assign read_data_reg_discontinue_lower = read_data_reg[TUSER_LOWER_OFFSET + 41];
   assign read_data_reg_tph_present_lower = read_data_reg[TUSER_LOWER_OFFSET + 42];  
   assign read_data_reg_tph_type_lower = read_data_reg[TUSER_LOWER_OFFSET + 44:
                                  TUSER_LOWER_OFFSET + 43];
   assign read_data_reg_tph_st_tag_lower = read_data_reg[TUSER_LOWER_OFFSET + 52:   
                                  TUSER_LOWER_OFFSET + 45];
  generate
    if (PARITY_ENABLE)
      begin
    assign read_data_reg_parity_lower = read_data_reg[TUSER_LOWER_OFFSET + 84:   
                                   TUSER_LOWER_OFFSET + 53];
    assign read_data_reg_eop_ptr_lower = read_data_reg[TUSER_LOWER_OFFSET + 87:
                                    TUSER_LOWER_OFFSET + 85];
      end
    else
      begin
    assign read_data_reg_parity_lower = 32'd0;
    assign read_data_reg_eop_ptr_lower = read_data_reg[TUSER_LOWER_OFFSET + 55:
                                    TUSER_LOWER_OFFSET + 53];
      end // else: !if(PARITY_ENABLE)
  endgenerate
      
   assign read_data_reg_first_be_upper = read_data_reg[TUSER_UPPER_OFFSET +3:
                               TUSER_UPPER_OFFSET];
   assign read_data_reg_last_be_upper = read_data_reg[TUSER_UPPER_OFFSET +7:
                              TUSER_UPPER_OFFSET +4];
   assign read_data_reg_byte_en_upper = read_data_reg[TUSER_UPPER_OFFSET +39:
                                 TUSER_UPPER_OFFSET +8];
   assign read_data_reg_sop_upper = read_data_reg[TUSER_UPPER_OFFSET + 40];
   assign read_data_reg_discontinue_upper = read_data_reg[TUSER_UPPER_OFFSET + 41];
   assign read_data_reg_tph_present_upper = read_data_reg[TUSER_UPPER_OFFSET + 42];  
   assign read_data_reg_tph_type_upper = read_data_reg[TUSER_UPPER_OFFSET + 44:
                                  TUSER_UPPER_OFFSET + 43];
   assign read_data_reg_tph_st_tag_upper = read_data_reg[TUSER_UPPER_OFFSET + 52:   
                                  TUSER_UPPER_OFFSET + 45];
  generate
    if (PARITY_ENABLE)
      begin
    assign read_data_reg_parity_upper = read_data_reg[TUSER_UPPER_OFFSET + 84:   
                                   TUSER_UPPER_OFFSET + 53];
    assign read_data_reg_eop_ptr_upper = read_data_reg[TUSER_UPPER_OFFSET + 87:
                               TUSER_UPPER_OFFSET + 85];
      end
    else
      begin
    assign read_data_reg_parity_upper = 32'd0;

    assign read_data_reg_eop_ptr_upper = read_data_reg[TUSER_UPPER_OFFSET + 55:
                               TUSER_UPPER_OFFSET + 53];
      end
  endgenerate

  generate
    if (PARITY_ENABLE)
      begin
    assign  read_data_reg_tlast_lower = read_data_reg[AXI4_CORE_DATA_WIDTH + AXI4_CORE_CQ_TKEEP_WIDTH +
                              AXI4_CORE_CQ_TUSER_WIDTH];
    assign     read_data_reg_tlast_upper = read_data_reg[AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_CQ_TKEEP_WIDTH*2 +
                              AXI4_CORE_CQ_TUSER_WIDTH*2 +2];
      end
    else
      begin
    assign  read_data_reg_tlast_lower = read_data_reg[AXI4_CORE_DATA_WIDTH + AXI4_CORE_CQ_TKEEP_WIDTH +
                              AXI4_CORE_CQ_TUSER_WIDTH -32];
    assign     read_data_reg_tlast_upper = read_data_reg[AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_CQ_TKEEP_WIDTH*2 +
                              AXI4_CORE_CQ_TUSER_WIDTH*2 +2 -64];
      end // else: !if(PARITY_ENABLE)
  endgenerate

   assign sop_in_lower_half = read_data_valid_reg[0] & read_data_reg_sop_lower;
   assign sop_in_upper_half = attr_straddle_en_i & read_data_valid_reg[1] & read_data_reg_sop_upper;

   assign eop_in_lower_half = read_data_valid_reg[0] & read_data_reg_tlast_lower;
   assign eop_in_upper_half = read_data_valid_reg[1] & read_data_reg_tlast_upper;
   
   assign read_data_out_first_be[3:0] = sop_in_lower_half? read_data_reg_first_be_lower: 
      sop_in_upper_half? read_data_reg_first_be_upper: 4'd0;
   assign read_data_out_first_be[7:4] = (sop_in_lower_half & sop_in_upper_half)?
      read_data_reg_first_be_upper: 4'd0;
   assign read_data_out_last_be[3:0] = sop_in_lower_half? read_data_reg_last_be_lower: 
      sop_in_upper_half? read_data_reg_last_be_upper: 4'd0;
   assign read_data_out_last_be[7:4] = (sop_in_lower_half & sop_in_upper_half)?
      read_data_reg_last_be_upper: 4'd0;
   assign read_data_out_byte_en[31:0] = read_data_valid_reg[0]? read_data_reg_byte_en_lower: 32'd0;
   assign read_data_out_byte_en[63:32] = read_data_valid_reg[1]? read_data_reg_byte_en_upper: 32'd0;
   
   assign read_data_out_is_sop[0] = sop_in_lower_half | sop_in_upper_half;
   assign read_data_out_is_sop[1] = sop_in_lower_half & sop_in_upper_half;

   assign read_data_out_is_sop0_ptr[1] = ~sop_in_lower_half & sop_in_upper_half;
   assign read_data_out_is_sop0_ptr[0] = 1'b0;
   assign read_data_out_is_sop1_ptr[1] = read_data_out_is_sop[1];
   assign read_data_out_is_sop1_ptr[0] = 1'b0;
   assign read_data_out_is_eop[0] = eop_in_lower_half | eop_in_upper_half;
   assign read_data_out_is_eop[1] = attr_straddle_en_i & eop_in_lower_half & eop_in_upper_half;
   assign read_data_out_is_eop0_ptr[3:0] = eop_in_lower_half? {1'b0, read_data_reg_eop_ptr_lower}:
      eop_in_upper_half? {1'b1, read_data_reg_eop_ptr_upper}: 4'd0;
   assign read_data_out_is_eop1_ptr[3:0] = (attr_straddle_en_i & eop_in_lower_half & eop_in_upper_half)?
      {1'b1, read_data_reg_eop_ptr_upper}: 4'd0;
   assign read_data_out_discontinue = (read_data_valid_reg[0] & read_data_reg_discontinue_lower) |
      (read_data_valid_reg[1] & read_data_reg_discontinue_upper);      

   assign read_data_out_tph_present[0] = sop_in_lower_half? read_data_reg_tph_present_lower:
      sop_in_upper_half? read_data_reg_tph_present_upper: 1'b0;
   assign read_data_out_tph_present[1] = (sop_in_lower_half & sop_in_upper_half)? read_data_reg_tph_present_upper: 1'b0;

   assign read_data_out_tph_type[1:0] = sop_in_lower_half? read_data_reg_tph_type_lower[1:0]:
      sop_in_upper_half? read_data_reg_tph_type_upper[1:0]: 2'd0;
   assign read_data_out_tph_type[3:2] = (sop_in_lower_half & sop_in_upper_half)? read_data_reg_tph_type_upper[1:0]: 2'd0;

   assign read_data_out_tph_st_tag[7:0] = sop_in_lower_half? read_data_reg_tph_st_tag_lower[7:0]:
      sop_in_upper_half? read_data_reg_tph_st_tag_upper[7:0]: 8'd0;
   assign read_data_out_tph_st_tag[15:8] = (sop_in_lower_half & sop_in_upper_half)? read_data_reg_tph_st_tag_upper[7:0]: 8'd0;

   assign read_data_out_parity[31:0] = read_data_valid_reg[0]? read_data_reg_parity_lower: 32'd0;
   assign read_data_out_parity[63:32] = read_data_valid_reg[1]? read_data_reg_parity_upper: 32'd0;

   assign read_data_out_tuser = {
                 read_data_out_parity[63:0],
                 read_data_out_tph_st_tag[15:0],
                 read_data_out_tph_type[3:0],
                 read_data_out_tph_present[1:0],
                 read_data_out_discontinue,
                 read_data_out_is_eop1_ptr[3:0],
                 read_data_out_is_eop0_ptr[3:0],
                 read_data_out_is_eop[1:0],
                 read_data_out_is_sop1_ptr[1:0],
                 read_data_out_is_sop0_ptr[1:0],
                 read_data_out_is_sop[1:0],
                 read_data_out_byte_en[63:0],
                 read_data_out_last_be[7:0],
                 read_data_out_first_be[7:0]
                 };


   assign read_data_out_tdata[AXI4_USER_DATA_WIDTH/2-1:0] = read_data_valid_reg[0]? read_data_reg[AXI4_CORE_DATA_WIDTH-1:0]:
      {AXI4_USER_DATA_WIDTH/2{1'b0}};
   assign read_data_out_tdata[AXI4_USER_DATA_WIDTH-1:AXI4_USER_DATA_WIDTH/2] = read_data_valid_reg[1]?
      read_data_reg[FIFO_READ_DATA_UPPER_OFFSET+AXI4_CORE_DATA_WIDTH-1:FIFO_READ_DATA_UPPER_OFFSET]: {AXI4_USER_DATA_WIDTH/2{1'b0}};
   
  assign  read_data_out_tkeep[AXI4_USER_CQ_TKEEP_WIDTH/2-1:0] = attr_straddle_en_i? {AXI4_USER_CQ_TKEEP_WIDTH/2{1'b1}}:
      read_data_valid_reg[0]? 
      read_data_reg[AXI4_CORE_DATA_WIDTH+AXI4_CORE_CQ_TKEEP_WIDTH-1:AXI4_CORE_DATA_WIDTH]: {AXI4_USER_CQ_TKEEP_WIDTH/2{1'b0}};
   assign read_data_out_tkeep[AXI4_USER_CQ_TKEEP_WIDTH-1:AXI4_USER_CQ_TKEEP_WIDTH/2] = attr_straddle_en_i? {AXI4_USER_CQ_TKEEP_WIDTH/2{1'b1}}:
      read_data_valid_reg[1]? 
      read_data_reg[FIFO_READ_TKEEP_UPPER_OFFSET+AXI4_CORE_CQ_TKEEP_WIDTH-1:FIFO_READ_TKEEP_UPPER_OFFSET]:
      {AXI4_USER_CQ_TKEEP_WIDTH/2{1'b0}};

   assign read_data_out_tlast = attr_straddle_en_i? 1'b0: (eop_in_lower_half | eop_in_upper_half);

   assign output_mux_in_data = {
                read_data_out_tlast,
                read_data_out_tuser,
                read_data_out_tkeep,
                read_data_out_tdata
                };

   // Instance of output MUX
   xp4_usp_smsw_512b_cq_output_mux #
     (
      .TCQ(TCQ),
      .IMPL_TARGET(IMPL_TARGET),
      .IN_DATA_WIDTH(OUTPUT_MUX_IN_DATA_WIDTH),
      .OUT_DATA_WIDTH(AXI4_USER_DATA_WIDTH),
      .TUSER_WIDTH(AXI4_USER_CQ_TUSER_WIDTH),
      .TKEEP_WIDTH(AXI4_USER_CQ_TKEEP_WIDTH)
      )
     pcie_4_0_512b_cq_output_mux_blk
       (
        .clk_i(user_clk_i),
        .reset_n_i(reset_n_user_clk_i),
        .link_down_reset_i(link_down_reset_i),
    .in_data_i(output_mux_in_data),
    .in_data_valid_i(read_data_valid_reg[0]),
        .attr_straddle_en_i(attr_straddle_en_i),

    .upstream_ready_o(output_mux_ready),
    .out_data_o(m_axis_cq_tdata_o),
        .out_data_valid_o(m_axis_cq_tvalid_o),
    .out_tuser_o(m_axis_cq_tuser_o),
    .out_tlast_o(m_axis_cq_tlast_o),
    .out_tkeep_o(m_axis_cq_tkeep_o),
    .downstream_ready_i(m_axis_cq_tready_i),
    
    .pcie_cq_np_req_i(pcie_cq_np_req_i),
    .pcie_cq_np_req_count_o(pcie_cq_np_req_count_o),
    .np_credit_received_o(cq_np_user_credit_rcvd_user_clk),
    .posted_req_delivered_o(posted_req_delivered_user_clk),
    .pipeline_empty_o(out_mux_pipeline_empty)
    );

   // Change clock domain for np_user_credit_rcvd signal
   always @(posedge user_clk2_i)
     if (~reset_n_user_clk2_i)
       cq_np_user_credit_rcvd_o <= #TCQ 1'b0;
     else
       if (user_clk_en_i)
     cq_np_user_credit_rcvd_o <= #TCQ cq_np_user_credit_rcvd_user_clk[0];
       else
     cq_np_user_credit_rcvd_o <= #TCQ cq_np_user_credit_rcvd_user_clk[1];

   // Change clock domain for posted_req_delivered signal
   always @(posedge user_clk2_i)
     if (~reset_n_user_clk2_i)
       posted_req_delivered_o <= #TCQ 1'b0;
     else
       if (user_clk_en_i)
     posted_req_delivered_o <= #TCQ posted_req_delivered_user_clk[0];
       else
     posted_req_delivered_o <= #TCQ posted_req_delivered_user_clk[1];

   assign pipeline_empty_user_clk = out_mux_pipeline_empty &&
      (read_data_valid_reg == 2'b00) &&
      ~fifo_read_data_valid &&
      ~fifo_in_data_valid_reg;

   always @(posedge user_clk2_i)
     if (~reset_n_user_clk2_i)
       pipeline_empty_core_clk <= #TCQ 1'b0;
     else
       pipeline_empty_core_clk <= #TCQ pipeline_empty_user_clk;

   always @(posedge user_clk2_i)
     if (~reset_n_user_clk2_i)
       cq_pipeline_empty_reg <= #TCQ 3'b111;
     else
       begin
      // Wait for pipeline empty signals to stay asserted for 3 cycles before signaling the output.
      cq_pipeline_empty_reg[0] <= #TCQ pipeline_empty_core_clk &
                      ~core_cq_tvalid_i &
                      ~core_cq_tvalid_reg_lower &
                      ~core_cq_tvalid_reg_upper;
         cq_pipeline_empty_reg[1] <= #TCQ cq_pipeline_empty_reg[0];
         cq_pipeline_empty_reg[2] <= #TCQ cq_pipeline_empty_reg[1];
      cq_pipeline_empty_o <= #TCQ &cq_pipeline_empty_reg;
       end // else: !if(~reset_n_user_clk2_i)
         

endmodule // pcie_4_0_512b_cq_intfc








   
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_512b_cq_output_mux.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_512b_cq_output_mux #(
   parameter TCQ = 100,
   parameter IMPL_TARGET = "SOFT",
   parameter IN_DATA_WIDTH = 512+183+16+1,    
   parameter OUT_DATA_WIDTH = 512,
   parameter TUSER_WIDTH = 183,
   parameter TKEEP_WIDTH = 16
   )
  (
    input  wire           clk_i // 250 MHz clock for client-facing interfaces
   ,input  wire           reset_n_i // Reset in the user clock domain
   ,input  wire           link_down_reset_i // Link went down

   ,input  wire           attr_straddle_en_i // Enable straddle

   ,input wire[IN_DATA_WIDTH-1:0] in_data_i
   ,input wire in_data_valid_i
   ,output wire upstream_ready_o

   ,output reg [OUT_DATA_WIDTH-1:0]  out_data_o
   ,output reg           out_data_valid_o
   ,output reg [TUSER_WIDTH-1:0] out_tuser_o
   ,output wire          out_tlast_o
   ,output wire [TKEEP_WIDTH-1:0] out_tkeep_o
   ,input  wire           downstream_ready_i

   ,input  wire [1:0]     pcie_cq_np_req_i // Client request to deliver NP TLP
   ,output reg [5:0]      pcie_cq_np_req_count_o // Current value of interface credit count for NP TLPs
   ,output reg [1:0]      np_credit_received_o // NP credit to TL
   ,output reg [1:0]      posted_req_delivered_o // Signals the delivery of a Posted Req on the CQ interface
   ,output wire           pipeline_empty_o // Indicates that the entire pipeline of the mux is empty
   );


   localparam MAX_CREDIT = 32;

   reg [1:0] output_fifo_occupancy;
   reg          output_fifo_write_ptr;
   reg          output_fifo_read_ptr;
   wire      output_fifo_full;
   wire      output_fifo_empty;

   reg [OUT_DATA_WIDTH-1:0] m_axis_cq_tdata_first_reg;
   reg [TKEEP_WIDTH-1:0]    m_axis_cq_tkeep_first_reg;
   reg [TUSER_WIDTH-1:0]    m_axis_cq_tuser_first_reg;
   reg                 m_axis_cq_tlast_first_reg;
   
   reg [OUT_DATA_WIDTH-1:0] m_axis_cq_tdata_second_reg;
   reg [TKEEP_WIDTH-1:0]    m_axis_cq_tkeep_second_reg;
   reg [TUSER_WIDTH-1:0]    m_axis_cq_tuser_second_reg;
   reg                 m_axis_cq_tlast_second_reg;
   
   wire             output_reg_mux_sel;

   wire [3:0]              output_reg_in_req_type0;
   wire [3:0]              output_reg_in_req_type1;
   
   wire              output_reg_in_req_type0_np;
   wire              output_reg_in_req_type1_np;

   wire              output_reg_in_sop0;
   wire              output_reg_in_sop1;
   wire              output_reg_in_eop0;
   wire              output_reg_in_eop1;
   wire              output_reg_in_error;

   reg [1:0]             pcie_cq_np_req_reg;
   reg                 tlp_in_progress;
   reg                 tlp_in_progress_type;

   reg [1:0]             np_tlp_count;
   
   wire [3:0]             out_req_type0;
   wire [3:0]             out_req_type1;
   reg                 m_axis_cq_tvalid_last;
   reg                 m_axis_cq_sop0_last;
   reg                 m_axis_cq_sop1_last;
   reg                 m_axis_cq_eop0_last;
   reg                 m_axis_cq_eop1_last;
   reg                 m_axis_cq_posted_type0_last;
   reg                 m_axis_cq_posted_type1_last;
   reg                 out_ready_reg;
   reg                 posted_tlp_in_progress;
   reg                 posted_tlp_in_progress_type;

  reg                 out_tlast_reg;
  reg [TKEEP_WIDTH-1:0]     out_tkeep_reg;

   //---------------------------------------------------------------------------------------------
   // Output FIFO
   // The main FIFO feeds into two read registers in the user clock domain, which are configured
   // as a 2-entry FIFO.
   // These are termed m_axis_cq_*_reg_first and m_axis_cq_*_reg_second.
   // These can be thought of as logical extensions of the main FIFO.
   //---------------------------------------------------------------------------------------------

   // Send signal to read from main FIFO into the output FIFO when the latter is not full.
   assign    upstream_ready_o = ~output_fifo_full;

   // Maintain write and read pointers
   always @(posedge clk_i)
     if (~reset_n_i)
       output_fifo_write_ptr <= #(TCQ) 1'b0;
     else if (link_down_reset_i)
       output_fifo_write_ptr <= #(TCQ) 1'b0;
     else
       if (in_data_valid_i & ~output_fifo_full)
	 output_fifo_write_ptr <= #(TCQ) ~output_fifo_write_ptr;

   always @(posedge clk_i)
     if (~reset_n_i)
       output_fifo_read_ptr <= #(TCQ) 1'b0;
     else if (link_down_reset_i)
       output_fifo_read_ptr <= #(TCQ) 1'b0;
     else
       if ((downstream_ready_i | ~out_data_valid_o) &
	   ~output_fifo_empty)
	 output_fifo_read_ptr <= #(TCQ) ~output_fifo_read_ptr;

    // Maintain FIFO occupancy
   always @(posedge clk_i)
     if (~reset_n_i)
       output_fifo_occupancy <= #(TCQ) 2'd0;
     else if (link_down_reset_i)
       output_fifo_occupancy <= #(TCQ) 2'd0;
     else
       if ((in_data_valid_i & ~output_fifo_full) &
       ~((downstream_ready_i | ~out_data_valid_o) &
         ~output_fifo_empty))
     output_fifo_occupancy <= #(TCQ) output_fifo_occupancy + 2'd1;
       else
     if (~(in_data_valid_i & ~output_fifo_full) &
         ((downstream_ready_i | ~out_data_valid_o) &
          ~output_fifo_empty))
       output_fifo_occupancy <= #(TCQ) output_fifo_occupancy - 2'd1;
   

   assign output_fifo_full = output_fifo_occupancy[1];
   assign output_fifo_empty = (output_fifo_occupancy == 2'b00);

   // Write data into the Output FIFO.                                                                                    
   always @(posedge clk_i)
     if (~reset_n_i)
       begin
          m_axis_cq_tdata_first_reg <= #(TCQ) {OUT_DATA_WIDTH{1'b0}};
          m_axis_cq_tdata_second_reg <= #(TCQ) {OUT_DATA_WIDTH{1'b0}};
          m_axis_cq_tkeep_first_reg <= #(TCQ) {TKEEP_WIDTH{1'b0}};
          m_axis_cq_tkeep_second_reg <= #(TCQ) {TKEEP_WIDTH{1'b0}};
          m_axis_cq_tuser_first_reg <= #(TCQ) {TUSER_WIDTH{1'b0}};
          m_axis_cq_tuser_second_reg <= #(TCQ) {TUSER_WIDTH{1'b0}};
          m_axis_cq_tlast_first_reg <= #(TCQ) 1'b0;
          m_axis_cq_tlast_second_reg <= #(TCQ) 1'b0;
       end
     else
        if (in_data_valid_i & ~output_fifo_full)
      begin
         case(output_fifo_write_ptr)
           1'b0:
         begin
            m_axis_cq_tdata_first_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH-1:0];
            m_axis_cq_tkeep_first_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH-1:OUT_DATA_WIDTH];
            m_axis_cq_tuser_first_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH+TUSER_WIDTH-1:OUT_DATA_WIDTH+TKEEP_WIDTH];
            m_axis_cq_tlast_first_reg <= #(TCQ) in_data_i[IN_DATA_WIDTH-1];
         end
           default:
         begin
            m_axis_cq_tdata_second_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH-1:0];
            m_axis_cq_tkeep_second_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH-1:OUT_DATA_WIDTH];
            m_axis_cq_tuser_second_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH+TUSER_WIDTH-1:OUT_DATA_WIDTH+TKEEP_WIDTH];
            m_axis_cq_tlast_second_reg <= #(TCQ) in_data_i[IN_DATA_WIDTH-1];
         end
         endcase // case(output_fifo_write_ptr)
      end // if (in_data_valid_i & ~output_fifo_full)
   
   // Output registers

   assign output_reg_mux_sel = output_fifo_read_ptr;

   always @(posedge clk_i)
     if (~reset_n_i)
       begin
      out_data_o <= #(TCQ) {OUT_DATA_WIDTH-1{1'b0}};
      out_tuser_o <= #(TCQ) {TUSER_WIDTH-1{1'b0}};
      out_tkeep_reg <= #(TCQ) {TKEEP_WIDTH-1{1'b0}};
      out_tlast_reg <= #(TCQ) 1'b0;
       end
     else
       if (~out_data_valid_o | downstream_ready_i)
     begin
        case(output_reg_mux_sel)
          1'b0:
        begin
           out_data_o <= #(TCQ) m_axis_cq_tdata_first_reg;
           out_tkeep_reg <= #(TCQ) m_axis_cq_tkeep_first_reg;
           out_tuser_o <= #(TCQ) m_axis_cq_tuser_first_reg;
           out_tlast_reg <= #(TCQ) m_axis_cq_tlast_first_reg;
        end
          default:
        begin
           out_data_o <= #(TCQ) m_axis_cq_tdata_second_reg;
           out_tkeep_reg <= #(TCQ) m_axis_cq_tkeep_second_reg;
           out_tuser_o <= #(TCQ) m_axis_cq_tuser_second_reg;
           out_tlast_reg <= #(TCQ) m_axis_cq_tlast_second_reg;
        end
        endcase // case(output_reg_mux_sel)
     end // if (~out_data_o | downstream_ready_i)

   always @(posedge clk_i)
     if (~reset_n_i)
       out_data_valid_o <= #(TCQ) 1'b0;
     else
       if (~out_data_valid_o | downstream_ready_i)
     out_data_valid_o <= #(TCQ) ~output_fifo_empty;

  assign out_tkeep_o =  attr_straddle_en_i? {TKEEP_WIDTH{1'b1}}: out_tkeep_reg;
  assign out_tlast_o =  attr_straddle_en_i? 1'b0: out_tlast_reg;

   //--------------------------------------------------------------------
   // NP credit management
   //-----------------------------------------------------------------------------------                

   // Decode packet Req Type as Posted/Non-Posted
   assign output_reg_in_req_type0 = in_data_i[78:75];
   assign output_reg_in_req_type1 = in_data_i[256+78:256+75];
   
   assign output_reg_in_req_type0_np = (output_reg_in_req_type0[3:0] != 4'd1) &&
	  (output_reg_in_req_type0[3:2] != 2'b11);
   assign output_reg_in_req_type1_np = (output_reg_in_req_type1[3:0] != 4'd1) &&
	  (output_reg_in_req_type1[3:2] != 2'b11);
  
   assign output_reg_in_sop0 = in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH+80];
   assign output_reg_in_sop1 = in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH+81];
   assign output_reg_in_eop0 = in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH+86];
   assign output_reg_in_eop1 = in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH+87];
   assign output_reg_in_error = in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH+95];  // discontinue  

   // Register the user input pcie_cq_np_req_i
   always @(posedge clk_i)
     if (~reset_n_i)
       pcie_cq_np_req_reg <= #(TCQ) 2'b00;
     else
       pcie_cq_np_req_reg <= #(TCQ) pcie_cq_np_req_i;

   // If a TLP is in progress from last beat, record its type.
  always @(posedge clk_i)
    if (~reset_n_i)
      begin
	tlp_in_progress <= 1'b0;
	tlp_in_progress_type <= 1'b0;
      end
  else if (in_data_valid_i & ~output_fifo_full)
    begin
      if (~tlp_in_progress)
	begin
	  if (output_reg_in_sop0 & ~output_reg_in_eop0)
            begin
              tlp_in_progress <= 1'b1;
              tlp_in_progress_type <= output_reg_in_req_type0_np;
            end
          else if (output_reg_in_sop1 & ~output_reg_in_eop1)
            begin
              tlp_in_progress <= 1'b1;
              tlp_in_progress_type <= output_reg_in_req_type1_np;
            end
          else
            begin
              tlp_in_progress <= 1'b0;
              tlp_in_progress_type <= 1'b0;
            end
	end // if (~tlp_in_progress)
      else
	begin
          if ((output_reg_in_eop0 & ~output_reg_in_sop0)|
	      output_reg_in_eop1)
	    tlp_in_progress <= 1'b0;
          if (output_reg_in_sop0)
	    tlp_in_progress_type <= output_reg_in_req_type1_np;
	end // else: !if(~tlp_in_progress)
    end // if (in_data_valid_i & ~output_fifo_full)
   
   // Determine number of NP TLPs being sent to user
   always @(*)
     begin
    case({output_reg_in_eop1, output_reg_in_eop0})
      2'd0: np_tlp_count = 2'd0;
      2'd1:
        begin
           if (~tlp_in_progress)
             begin
               if (output_reg_in_req_type0_np & ~output_reg_in_error)
		 np_tlp_count = 2'd1;
               else
		 np_tlp_count = 2'd0;
             end
           else
             begin
               if (tlp_in_progress_type & ~output_reg_in_error)
		 np_tlp_count = 2'd1;
               else
		 np_tlp_count = 2'd0;
             end // else: !if(~tlp_in_progress)
	end // case: 2'd1
      
      default: //2'd3
        begin
           if (~tlp_in_progress)
             begin
               if (output_reg_in_req_type0_np & output_reg_in_req_type1_np)
		 np_tlp_count = 2'd2;
               else if (output_reg_in_req_type0_np | output_reg_in_req_type1_np)
		 np_tlp_count = 2'd1;
               else
		 np_tlp_count = 2'd0;
             end
           else
             begin
               if (tlp_in_progress_type & output_reg_in_req_type1_np)
		 np_tlp_count = 2'd2;
               else if (tlp_in_progress_type | output_reg_in_req_type1_np)
		 np_tlp_count = 2'd1;
               else
		 np_tlp_count = 2'd0;
             end // else: !if(~tlp_in_progress)
        end // case: default
    endcase // case({output_reg_in_eop1, output_reg_in_eop0})
     end // always @ (*)

   // Maintain current NP credit
   always @(posedge clk_i)
     if (~reset_n_i)
       begin
      pcie_cq_np_req_count_o <= 6'd0;
       end
     else if (link_down_reset_i)
       begin
      pcie_cq_np_req_count_o <= 6'd0;
       end
     else
       if (in_data_valid_i & ~output_fifo_full)
     begin
        casez({np_tlp_count, pcie_cq_np_req_reg})
          4'b00_01:
        begin
           // No TLPs being delivered, user provided 1 credit
           if (pcie_cq_np_req_count_o != MAX_CREDIT[5:0])
             pcie_cq_np_req_count_o <= pcie_cq_np_req_count_o + 6'd1;
        end
          4'b00_1?:
        begin
           // No TLPs being delivered, user provided 2 credits
           if (pcie_cq_np_req_count_o <= (MAX_CREDIT-2))
             pcie_cq_np_req_count_o <= pcie_cq_np_req_count_o + 6'd2;
           else
             pcie_cq_np_req_count_o <= MAX_CREDIT[5:0];
        end
          4'b01_00:
        begin
           // One NP TLP being delivered, user provided no credit
           if (pcie_cq_np_req_count_o != 6'd0)
             pcie_cq_np_req_count_o <= pcie_cq_np_req_count_o - 6'd1;
        end
          4'b01_1?:
        begin
           // One NP TLP being delivered, user provided 2 credits
           if (pcie_cq_np_req_count_o != MAX_CREDIT[5:0])
             pcie_cq_np_req_count_o <= pcie_cq_np_req_count_o + 6'd1;
        end
          4'b1?_00:
        begin
           // Two NP TLP being delivered, user provided no credit.
           // Decrement by 2.
           if (pcie_cq_np_req_count_o[5:1] != 5'd0)
             pcie_cq_np_req_count_o <= pcie_cq_np_req_count_o - 6'd2;
           else
             pcie_cq_np_req_count_o[0] <= 1'b0;
        end          
          4'b1?_01:
        begin
           // Two NP TLP being delivered, user provided 1 credit.
           // Decrement by 1.
           if (pcie_cq_np_req_count_o != 6'd0)
             pcie_cq_np_req_count_o <= pcie_cq_np_req_count_o - 6'd1;
        end
        endcase // casez({np_tlp_count, pcie_cq_np_req_reg})
     end // if (in_data_valid_i & ~output_fifo_full)
       else
     begin
       casez(pcie_cq_np_req_reg)
         2'b01:
           begin
         // No TLPs being delivered, user provided 1 credit
         if (pcie_cq_np_req_count_o != MAX_CREDIT[5:0])
           pcie_cq_np_req_count_o <= pcie_cq_np_req_count_o + 6'd1;
           end
         2'b1?:
           begin
         // No TLPs being delivered, user provided 2 credits
         if (pcie_cq_np_req_count_o <= (MAX_CREDIT-2))
           pcie_cq_np_req_count_o <= pcie_cq_np_req_count_o + 6'd2;
         else
           pcie_cq_np_req_count_o <= MAX_CREDIT[5:0];
           end
         default:
           begin
           end
       endcase // casez(pcie_cq_np_req_reg)
     end // else: !if(in_data_valid_i & ~output_fifo_full)

  // Send indication to Transaction Layer when user issues more credit
   always @(posedge clk_i)
     if (~reset_n_i)
       np_credit_received_o <= 2'b00;
     else
       if (in_data_valid_i & ~output_fifo_full)
     begin
        casez({np_tlp_count, pcie_cq_np_req_reg})
          4'b00_01:
        // No TLPs being delivered, user provided 1 credit
        begin
           // Provide credit to TL when credit count has not saturated
           if (pcie_cq_np_req_count_o == MAX_CREDIT[5:0])
             np_credit_received_o <= 2'b00;
           else
             np_credit_received_o <= 2'b01;
        end
          4'b00_1?:
        // No TLPs being delivered, user provided 2 credits
        begin
           // Provide credit to TL when credit count has not saturated
           if (pcie_cq_np_req_count_o == MAX_CREDIT[5:0])
             np_credit_received_o <= 2'b00;
           else if (pcie_cq_np_req_count_o == (MAX_CREDIT -1))
             // Provide 1 credit.
             np_credit_received_o <= 2'b01;
           else
             // Provide 2 credits.
             np_credit_received_o <= 2'b11;
        end // case: 4'b00_1x
          4'b01_01:
        // 1 TLP being delivered, user provided 1 credit
        begin
           // Always provide 1 credit to TL
           np_credit_received_o <= 2'b01;
        end
          4'b01_1?:
        // 1 TLP being delivered, user provided 2 credits
        begin
           // Provide 1 credit to TL when credit count has not saturated
           if (pcie_cq_np_req_count_o == MAX_CREDIT[5:0])
             np_credit_received_o <= 2'b01;
           else
             np_credit_received_o <= 2'b11;
        end
          4'b1?_01:
        // 2 TLPs being delivered, user provided 1 credit
        begin
           // Always provide 1 credit to TL
           np_credit_received_o <= 2'b01;
        end
          4'b1?_1?:
        // 2 TLPs being delivered, user provided 2 credits
        begin
           // Always provide 2 credits to TL
           np_credit_received_o <= 2'b11;
        end
          default:
        begin
           np_credit_received_o <= 2'b00;
        end
        endcase // casez({np_tlp_count, pcie_cq_np_req_reg})
     end // if (in_data_valid_i & ~output_fifo_full)
       else
     begin
       casez(pcie_cq_np_req_reg)
         2'b01:
           begin
         // No TLPs being delivered, user provided 1 credit
         if (pcie_cq_np_req_count_o != MAX_CREDIT[5:0])
           np_credit_received_o <= 2'b01;
         else
           np_credit_received_o <= 2'b00;
           end
         2'b1?:
           begin
         // No TLPs being delivered, user provided 2 credits.
         // Provide credit to TL when credit count has not saturated
         if (pcie_cq_np_req_count_o == MAX_CREDIT[5:0])
           np_credit_received_o <= 2'b00;
         else if (pcie_cq_np_req_count_o == (MAX_CREDIT -1))
           // Provide 1 credit.
           np_credit_received_o <= 2'b01;
         else
           // Provide 2 credits.
           np_credit_received_o <= 2'b11;
           end // case: 4'b00_1?
         default:
           begin
         np_credit_received_o <= 2'b00;
           end
       endcase // casez(pcie_cq_np_req_reg)
     end // else: !if(in_data_valid_i & ~output_fifo_full)

 //-------------------------------------------------------------------------------------------
   // Generate indication when a Posted request is delivered to the user

   assign out_req_type0 = out_data_o[78:75];
   assign out_req_type1 = out_data_o[256+78:256+75];

   always @(posedge clk_i)
     if (~reset_n_i)
       begin
      m_axis_cq_tvalid_last <= 1'b0;
      m_axis_cq_sop0_last <= 1'b0;
      m_axis_cq_sop1_last <= 1'b0;
      m_axis_cq_eop0_last <= 1'b0;
      m_axis_cq_eop1_last <= 1'b0;
      m_axis_cq_posted_type0_last <= 1'b0;
      m_axis_cq_posted_type1_last <= 1'b0;
       end
     else
       begin
      m_axis_cq_tvalid_last <= out_data_valid_o;
      m_axis_cq_sop0_last <= out_tuser_o[80];
      m_axis_cq_sop1_last <= out_tuser_o[81];
      m_axis_cq_eop0_last <= out_tuser_o[86];
      m_axis_cq_eop1_last <= out_tuser_o[87];
      m_axis_cq_posted_type0_last <= (out_req_type0[3:0] == 4'd1) || (out_req_type0[3:2] == 2'b11);
      m_axis_cq_posted_type1_last <= (out_req_type1[3:0] == 4'd1) || (out_req_type1[3:2] == 2'b11);
       end // else: !if(~reset_n_i)

   // Register ready
   always @(posedge clk_i)
     if (~reset_n_i)
       out_ready_reg <= 1'b0;
     else
       out_ready_reg <= downstream_ready_i;

   always @(posedge clk_i)
     if (~reset_n_i)
       begin
      posted_tlp_in_progress <= 1'b0;
      posted_tlp_in_progress_type <= 1'b0;
       end
     else if (link_down_reset_i)
       posted_tlp_in_progress <= 1'b0;
     else if (m_axis_cq_tvalid_last & out_ready_reg)
       begin
          if (~posted_tlp_in_progress)
        begin
           if (m_axis_cq_sop0_last & ~m_axis_cq_eop0_last)
         begin
            posted_tlp_in_progress <= 1'b1;
            posted_tlp_in_progress_type <=  m_axis_cq_posted_type0_last;
         end
           else if (m_axis_cq_sop1_last & ~m_axis_cq_eop1_last)
         begin
            posted_tlp_in_progress <= 1'b1;
            posted_tlp_in_progress_type <=  m_axis_cq_posted_type1_last;
         end
           else
         posted_tlp_in_progress <= 1'b0;
        end // if (~posted_tlp_in_progress)
      else
        begin
           if ((m_axis_cq_eop0_last & ~m_axis_cq_sop0_last) |
           m_axis_cq_eop1_last)
         posted_tlp_in_progress <= 1'b0;

           if (m_axis_cq_sop0_last)
         posted_tlp_in_progress_type <= m_axis_cq_posted_type1_last;
        end // else: !if(~posted_tlp_in_progress)
       end // if (m_axis_cq_tvalid_last & out_ready_reg)

   always @(posedge clk_i)
     if (~reset_n_i)
       posted_req_delivered_o <= 2'b00;
     else if (m_axis_cq_tvalid_last & out_ready_reg)
       begin
          if (~posted_tlp_in_progress)
        begin
          if ((m_axis_cq_sop0_last & m_axis_cq_posted_type0_last & m_axis_cq_eop0_last) &
          (m_axis_cq_sop1_last & m_axis_cq_posted_type1_last & m_axis_cq_eop1_last))
        // Two Complete TLPs in this beat.
        posted_req_delivered_o <= 2'b11;
          else if ((m_axis_cq_sop0_last & m_axis_cq_posted_type0_last & m_axis_cq_eop0_last) |
               (m_axis_cq_sop1_last & m_axis_cq_posted_type1_last & m_axis_cq_eop1_last))
        // Single TLP beginning and ending in this beat.
        posted_req_delivered_o <= 2'b01;
          else
        // No Posted TLP ending in this beat
        posted_req_delivered_o <= 2'b00;
        end // if (~tlp_in_progress)
      else
        begin
               if ((posted_tlp_in_progress_type & m_axis_cq_eop0_last) &
           (m_axis_cq_sop0_last & m_axis_cq_posted_type1_last & m_axis_cq_eop1_last))
         // TLP in progress ended in this cycle, and a new TLP started and ended.
         posted_req_delivered_o <= 2'b11;
               else if ((posted_tlp_in_progress_type & m_axis_cq_eop0_last) |
            (m_axis_cq_sop0_last & m_axis_cq_posted_type1_last & m_axis_cq_eop1_last))
         posted_req_delivered_o <= 2'b01;
           else
         posted_req_delivered_o <= 2'b00;
        end // else: !if(~posted_tlp_in_progress)
       end // if (m_axis_cq_tvalid_last & out_ready_reg)
     else
       posted_req_delivered_o <= 2'b00;

  assign pipeline_empty_o = output_fifo_empty && ~out_data_valid_o && ~m_axis_cq_tvalid_last && (posted_req_delivered_o == 2'b00);


endmodule // pcie_4_0_512b_cq_output_mux
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_512b_rc_intfc.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_512b_rc_intfc #(
   parameter TCQ = 100,
   parameter IMPL_TARGET = "SOFT",
   parameter AXISTEN_IF_EXT_512_INTFC_RAM_STYLE = "SRL",
   parameter AXI4_USER_DATA_WIDTH = 512,
   parameter AXI4_CORE_DATA_WIDTH = 256,
   parameter AXI4_USER_RC_TUSER_WIDTH = 161,                
   parameter AXI4_CORE_RC_TUSER_WIDTH = 75,
   parameter AXI4_USER_RC_TKEEP_WIDTH = 16,
   parameter AXI4_CORE_RC_TKEEP_WIDTH = 8,                
   parameter AXI4_CORE_RC_TREADY_WIDTH = 22,
   parameter PARITY_ENABLE = 0                
     ) 
  (
    input  wire           user_clk2_i // 500 MHz clock for core-facing interfaces
   ,input  wire           user_clk_i // 250 MHz clock for client-facing interfaces
   ,input  wire           user_clk_en_i // User clock enable for clock domain crossing
   ,input  wire           reset_n_user_clk_i // Reset in the user clock domain
   ,input  wire           reset_n_user_clk2_i // Reset in the user clock2 domain
   ,input  wire           link_down_reset_i // Link went down
   // Attributes
   ,input  wire           attr_straddle_en_i // Enable straddle
   ,input  wire           attr_4tlp_straddle_en_i  // Enable 4-tlp straddle
   ,input wire [1:0]      attr_alignment_mode_i // Payload alignment mode
                                                // (00= Dword-aligned, 10 = 128b address-aligned)
   //-----------------------------------------------------------------------------------------------
   // Client-side signals
   //-----------------------------------------------------------------------------------------------
   ,output wire [511:0]   m_axis_rc_tdata_o
   ,output wire           m_axis_rc_tvalid_o
   ,output wire [160:0]   m_axis_rc_tuser_o
   ,output wire           m_axis_rc_tlast_o
   ,output wire [15:0]    m_axis_rc_tkeep_o
   ,input  wire           m_axis_rc_tready_i
   //-----------------------------------------------------------------------------------------------
   // Core-side signals
   //-----------------------------------------------------------------------------------------------
   ,input  wire [255:0]   core_rc_tdata_i
   ,input  wire           core_rc_tvalid_i
   ,input  wire [74:0]    core_rc_tuser_i
   ,input  wire           core_rc_tlast_i
   ,input  wire [7:0]     core_rc_tkeep_i
   ,output wire [21:0]     core_rc_tready_o
   // Completion delivered indications
   ,output reg [1:0]      compl_delivered_o // Completions delivered to user
                                            // 00 = No Compl, 01 = 1 Compl, 11 = 2 Completions
   ,output reg [7:0]      compl_delivered_tag0_o// Tag associated with first delivered Completion
   ,output reg [7:0]      compl_delivered_tag1_o// Tag associated with second delivered Completion
   );

   localparam FIFO_WIDTH = PARITY_ENABLE? (AXI4_CORE_DATA_WIDTH + (AXI4_CORE_RC_TUSER_WIDTH+1) +
                       AXI4_CORE_RC_TKEEP_WIDTH + 1)*2 +2 :
               (AXI4_CORE_DATA_WIDTH + (AXI4_CORE_RC_TUSER_WIDTH+1) + 
                AXI4_CORE_RC_TKEEP_WIDTH + 1)*2 +2 -64;

   localparam TUSER_LOWER_OFFSET = AXI4_CORE_DATA_WIDTH + AXI4_CORE_RC_TKEEP_WIDTH;
   localparam TUSER_UPPER_OFFSET = PARITY_ENABLE? AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_RC_TKEEP_WIDTH*2 +
                   (AXI4_CORE_RC_TUSER_WIDTH+1) +2:
                   AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_RC_TKEEP_WIDTH*2 +
                   (AXI4_CORE_RC_TUSER_WIDTH+1) +2 -32;
   
  localparam FIFO_READ_DATA_UPPER_OFFSET = PARITY_ENABLE?
                   AXI4_CORE_DATA_WIDTH + AXI4_CORE_RC_TKEEP_WIDTH + (AXI4_CORE_RC_TUSER_WIDTH+1) +2:
                   AXI4_CORE_DATA_WIDTH + AXI4_CORE_RC_TKEEP_WIDTH + (AXI4_CORE_RC_TUSER_WIDTH+1) +2 -32;
  
  localparam FIFO_READ_TKEEP_UPPER_OFFSET = PARITY_ENABLE?
                    AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_RC_TKEEP_WIDTH + (AXI4_CORE_RC_TUSER_WIDTH+1) +2:
                                    AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_RC_TKEEP_WIDTH + (AXI4_CORE_RC_TUSER_WIDTH+1) +2 -32;

   localparam OUTPUT_MUX_IN_DATA_WIDTH = AXI4_USER_DATA_WIDTH +
                     AXI4_USER_RC_TKEEP_WIDTH +
                     AXI4_USER_RC_TUSER_WIDTH + 1;


   (* KEEP = "true" *) reg [AXI4_CORE_RC_TREADY_WIDTH-1:0] core_rc_tready_reg;
   (* KEEP = "true" *) reg core_rc_tready_user_clk2;

   reg [AXI4_CORE_DATA_WIDTH-1:0] core_rc_tdata_reg_upper;
   reg [AXI4_CORE_DATA_WIDTH-1:0] core_rc_tdata_reg_lower;
   reg [AXI4_CORE_RC_TUSER_WIDTH-1:0] core_rc_tuser_reg_upper;
   reg [AXI4_CORE_RC_TUSER_WIDTH-1:0] core_rc_tuser_reg_lower;
   reg                       core_rc_tlast_reg_upper;
   reg                       core_rc_tlast_reg_lower;
   reg [AXI4_CORE_RC_TKEEP_WIDTH-1:0] core_rc_tkeep_reg_upper;
   reg [AXI4_CORE_RC_TKEEP_WIDTH-1:0] core_rc_tkeep_reg_lower;
   reg                       core_rc_tvalid_reg_upper;
   reg                       core_rc_tvalid_reg_lower;

   reg [AXI4_CORE_DATA_WIDTH-1:0] core_rc_tdata_reg_upper_user_clk;
   reg [AXI4_CORE_DATA_WIDTH-1:0] core_rc_tdata_reg_lower_user_clk;
   reg [AXI4_CORE_RC_TUSER_WIDTH-1:0] core_rc_tuser_reg_upper_user_clk;
   reg [AXI4_CORE_RC_TUSER_WIDTH-1:0] core_rc_tuser_reg_lower_user_clk;
   reg                       core_rc_tlast_reg_upper_user_clk;
   reg                       core_rc_tlast_reg_lower_user_clk;
   reg [AXI4_CORE_RC_TKEEP_WIDTH-1:0] core_rc_tkeep_reg_upper_user_clk;
   reg [AXI4_CORE_RC_TKEEP_WIDTH-1:0] core_rc_tkeep_reg_lower_user_clk;
   reg                       core_rc_tvalid_reg_upper_user_clk;
   reg                       core_rc_tvalid_reg_lower_user_clk;
   wire [2:0]                core_rc_eop_ptr_upper;
   wire [2:0]                core_rc_eop_ptr_lower;
   wire [AXI4_CORE_RC_TUSER_WIDTH-1:0] core_rc_tuser_reg_upper_user_clk_int;
   wire [AXI4_CORE_RC_TUSER_WIDTH-1:0] core_rc_tuser_reg_lower_user_clk_int;


   wire                   fifo_almost_full_user_clk;

  reg                       core_rc_pkt_in_progress;
  wire                       core_rc_pkt_in_progress_upper;
  wire                       core_rc_tuser_sop0_lower;
  wire                       core_rc_tuser_sop1_lower;
  wire                       core_rc_tuser_eop0_lower;
  wire                       core_rc_tuser_eop1_lower;
  wire                       core_rc_tuser_sop0_upper;
  wire                       core_rc_tuser_sop1_upper;
  wire                       core_rc_tuser_eop0_upper;
  wire                       core_rc_tuser_eop1_upper;
  
  wire                       core_rc_tuser_reg_sop0_ptr_lower;
  wire                       core_rc_tuser_reg_sop0_ptr_upper;

   wire [FIFO_WIDTH-1:0]           fifo_in_data;
   reg                       fifo_in_data_valid;
   reg                       fifo_read_en;
   wire                   fifo_read_data_valid;
   wire [FIFO_WIDTH-1:0]           fifo_read_data;

   wire                   read_sop0_lower;
   wire                    read_sop0_ptr_lower;
   wire                   read_sop1_lower;
   wire                   read_discontinue_lower;
   wire                    read_eop0_lower;
   wire                    read_eop1_lower;
   wire                    read_eop_lower;
   wire                   read_tlast_lower;
   wire                   read_tlast_upper;
   wire                   read_data_valid_lower;
   wire                   read_data_valid_upper;

   wire                   read_sop0_upper;
   wire                    read_sop0_ptr_upper;
   wire                   read_sop1_upper;
   wire                   read_sop_upper;
   wire                   read_discontinue_upper;
   wire                    read_eop0_upper;
   wire                    read_eop1_upper;
   wire                    read_eop_upper;

   reg [1:0]                   read_data_valid_reg;
   reg [FIFO_WIDTH-1:0]           read_data_reg;
   reg [FIFO_WIDTH/2-1:0]           saved_data_reg;
   reg                       saved_eop;
   reg                       saved_err;
   
   wire [31:0]                   read_data_reg_byte_en_lower;
   wire                    read_data_reg_sop0_lower;
   wire                    read_data_reg_sop0_ptr_lower;
   wire                    read_data_reg_sop1_lower;
   wire                    read_data_reg_discontinue_lower;
   wire [31:0]                   read_data_reg_parity_lower;
   wire                    read_data_reg_eop0_lower;
   wire [2:0]                   read_data_reg_eop0_ptr_lower;
   wire                    read_data_reg_eop1_lower;
   wire [2:0]                   read_data_reg_eop1_ptr_lower;

   wire [31:0]                   read_data_reg_byte_en_upper;
   wire                    read_data_reg_sop0_upper;
   wire                    read_data_reg_sop0_ptr_upper;
   wire                    read_data_reg_sop1_upper;
   wire                    read_data_reg_discontinue_upper;
   wire [31:0]                   read_data_reg_parity_upper;
   wire                    read_data_reg_eop0_upper;
   wire [2:0]                   read_data_reg_eop0_ptr_upper;
   wire                    read_data_reg_eop1_upper;
   wire [2:0]                   read_data_reg_eop1_ptr_upper;

  wire                       read_data_reg_tlast_lower;
  wire                       read_data_reg_tlast_upper;

   wire [63:0]                   read_data_out_byte_en;
   wire [3:0]                   read_data_out_is_sop;
   wire [1:0]                   read_data_out_is_sop0_ptr;
   wire [1:0]                   read_data_out_is_sop1_ptr;
   wire [1:0]                   read_data_out_is_sop2_ptr;
   wire [1:0]                   read_data_out_is_sop3_ptr;
   wire [3:0]                   read_data_out_is_eop;
   wire [3:0]                   read_data_out_is_eop0_ptr;
   wire [3:0]                   read_data_out_is_eop1_ptr;
   wire [3:0]                   read_data_out_is_eop2_ptr;
   wire [3:0]                   read_data_out_is_eop3_ptr;
   wire                   read_data_out_discontinue;
   wire [63:0]                   read_data_out_parity;
   
   wire [ AXI4_USER_RC_TUSER_WIDTH-1:0] read_data_out_tuser;
   wire [ AXI4_USER_DATA_WIDTH-1:0]     read_data_out_tdata;
   wire [ AXI4_USER_RC_TKEEP_WIDTH-1:0] read_data_out_tkeep;
   wire                 read_data_out_tlast;
   
   wire [OUTPUT_MUX_IN_DATA_WIDTH-1:0]     output_mux_in_data;

   wire                 output_mux_ready;
   
  wire [3:0]                 pcie_compl_delivered_user_clk;
  wire [7:0]                 pcie_compl_delivered_tag0_user_clk;
  wire [7:0]                 pcie_compl_delivered_tag1_user_clk;
  wire [7:0]                 pcie_compl_delivered_tag2_user_clk;
  wire [7:0]                 pcie_compl_delivered_tag3_user_clk;

   // Read State Machine states
   localparam                           IDLE = 2'd0;
   localparam                           EXPECT_NEW_WORD = 2'd1;
   localparam                           SEND_SAVED_HALF_WORD = 2'd2;
   localparam                           WAIT_FOR_UPPER_HALF = 2'd3;
   reg [1:0]                 read_state;

   // Capture incoming data from core at 500 MHz into upper and lower registers
   always @(posedge user_clk2_i)
     if (~reset_n_user_clk2_i)
       begin
      core_rc_tdata_reg_upper <= #TCQ {AXI4_CORE_DATA_WIDTH{1'b0}};
      core_rc_tdata_reg_lower <= #TCQ {AXI4_CORE_DATA_WIDTH{1'b0}};
      core_rc_tuser_reg_upper <= #TCQ {AXI4_CORE_RC_TUSER_WIDTH{1'b0}};
      core_rc_tuser_reg_lower <= #TCQ {AXI4_CORE_RC_TUSER_WIDTH{1'b0}};
      core_rc_tkeep_reg_upper <= #TCQ {AXI4_CORE_RC_TKEEP_WIDTH{1'b0}};
      core_rc_tkeep_reg_lower <= #TCQ {AXI4_CORE_RC_TKEEP_WIDTH{1'b0}};
      core_rc_tlast_reg_upper <= #TCQ 1'b0;
      core_rc_tlast_reg_lower <= #TCQ 1'b0;
       core_rc_tvalid_reg_upper <= #TCQ 1'b0;
      core_rc_tvalid_reg_lower <= #TCQ 1'b0;
       end // if (~reset_n_user_clk_i)
     else
       if (user_clk_en_i)
     begin
        core_rc_tdata_reg_lower <= #TCQ core_rc_tdata_i;
        core_rc_tuser_reg_lower <= #TCQ core_rc_tuser_i;
        core_rc_tkeep_reg_lower <= #TCQ core_rc_tkeep_i;
        core_rc_tlast_reg_lower <= #TCQ core_rc_tlast_i;
        core_rc_tvalid_reg_lower <= #TCQ core_rc_tvalid_i & core_rc_tready_user_clk2;
     end
       else
     begin
        core_rc_tdata_reg_upper <= #TCQ core_rc_tdata_i;
        core_rc_tuser_reg_upper <= #TCQ core_rc_tuser_i;
        core_rc_tkeep_reg_upper <= #TCQ core_rc_tkeep_i;
        core_rc_tlast_reg_upper <= #TCQ core_rc_tlast_i;
        core_rc_tvalid_reg_upper <= #TCQ core_rc_tvalid_i & core_rc_tready_user_clk2;
     end // else: !if(user_clk_en_i)

  // Transfer to 250 MHz user_clk domain
     always @(posedge user_clk_i)
     if (~reset_n_user_clk_i)
       begin
     core_rc_tdata_reg_upper_user_clk <= #TCQ {AXI4_CORE_DATA_WIDTH{1'b0}};
     core_rc_tdata_reg_lower_user_clk <= #TCQ {AXI4_CORE_DATA_WIDTH{1'b0}};
     core_rc_tuser_reg_upper_user_clk <= #TCQ {AXI4_CORE_RC_TUSER_WIDTH{1'b0}};
     core_rc_tuser_reg_lower_user_clk <= #TCQ {AXI4_CORE_RC_TUSER_WIDTH{1'b0}};
     core_rc_tkeep_reg_upper_user_clk <= #TCQ {AXI4_CORE_RC_TKEEP_WIDTH{1'b0}};
     core_rc_tkeep_reg_lower_user_clk <= #TCQ {AXI4_CORE_RC_TKEEP_WIDTH{1'b0}};
     core_rc_tlast_reg_upper_user_clk <= #TCQ 1'b0;
     core_rc_tlast_reg_lower_user_clk <= #TCQ 1'b0;
      core_rc_tvalid_reg_upper_user_clk <= #TCQ 1'b0;
     core_rc_tvalid_reg_lower_user_clk <= #TCQ 1'b0;
     fifo_in_data_valid <= #TCQ 1'b0;
       end // if (~reset_n_user_clk_i)
     else
       begin
            core_rc_tdata_reg_upper_user_clk <= #TCQ core_rc_tdata_reg_upper;
     core_rc_tdata_reg_lower_user_clk <= #TCQ core_rc_tdata_reg_lower;
     core_rc_tuser_reg_upper_user_clk <= #TCQ core_rc_tuser_reg_upper;
     core_rc_tuser_reg_lower_user_clk <= #TCQ core_rc_tuser_reg_lower;
     core_rc_tkeep_reg_upper_user_clk <= #TCQ core_rc_tkeep_reg_upper;
     core_rc_tkeep_reg_lower_user_clk <= #TCQ core_rc_tkeep_reg_lower;
     core_rc_tlast_reg_upper_user_clk <= #TCQ core_rc_tlast_reg_upper;
     core_rc_tlast_reg_lower_user_clk <= #TCQ core_rc_tlast_reg_lower;
      core_rc_tvalid_reg_upper_user_clk <= #TCQ core_rc_tvalid_reg_upper;
     core_rc_tvalid_reg_lower_user_clk <= #TCQ core_rc_tvalid_reg_lower;
     fifo_in_data_valid <= #TCQ core_rc_tvalid_reg_upper | core_rc_tvalid_reg_lower;
       end // else: !if(~reset_n_user_clk_i)
  
  assign core_rc_eop_ptr_lower   = (core_rc_tkeep_reg_lower_user_clk[7])? 3'd7:
                                   (core_rc_tkeep_reg_lower_user_clk[6])? 3'd6:
                                   (core_rc_tkeep_reg_lower_user_clk[5])? 3'd5:
                                   (core_rc_tkeep_reg_lower_user_clk[4])? 3'd4:
                                   (core_rc_tkeep_reg_lower_user_clk[3])? 3'd3:
                                   (core_rc_tkeep_reg_lower_user_clk[2])? 3'd2:
                                   (core_rc_tkeep_reg_lower_user_clk[1])? 3'd1: 3'd0;
  assign core_rc_eop_ptr_upper   = (core_rc_tkeep_reg_upper_user_clk[7])? 3'd7:
                                   (core_rc_tkeep_reg_upper_user_clk[6])? 3'd6:
                                   (core_rc_tkeep_reg_upper_user_clk[5])? 3'd5:
                                   (core_rc_tkeep_reg_upper_user_clk[4])? 3'd4:
                                   (core_rc_tkeep_reg_upper_user_clk[3])? 3'd3:
                                   (core_rc_tkeep_reg_upper_user_clk[2])? 3'd2:
                                   (core_rc_tkeep_reg_upper_user_clk[1])? 3'd1: 3'd0;
  assign core_rc_tuser_reg_lower_user_clk_int   = (~attr_4tlp_straddle_en_i)? {core_rc_tuser_reg_lower_user_clk[AXI4_CORE_RC_TUSER_WIDTH-1:42],
                                                                               4'd0,   // [41:38], is_eop_1[3:0]
                                                                               core_rc_eop_ptr_lower, // [37:35]
                                                                               core_rc_tlast_reg_lower_user_clk,  // [34]
                                                                               1'b0,   // [33], is_sop_1
                                                                               core_rc_tuser_reg_lower_user_clk[32:0]}:
                                                                              core_rc_tuser_reg_lower_user_clk;
  assign core_rc_tuser_reg_upper_user_clk_int   = (~attr_4tlp_straddle_en_i)? {core_rc_tuser_reg_upper_user_clk[AXI4_CORE_RC_TUSER_WIDTH-1:42],
                                                                               4'd0,   // [41:38], is_eop_1[3:0]
                                                                               core_rc_eop_ptr_upper, // [37:35]
                                                                               core_rc_tlast_reg_upper_user_clk,  // [34]
                                                                               1'b0,   // [33], is_sop_1
                                                                               core_rc_tuser_reg_upper_user_clk[32:0]}:
                                                                              core_rc_tuser_reg_upper_user_clk;
  // Generate SOP0 Pointer for lower and upper halves.
  // This requires keeping track of whether a packet is continuing from the last beat.
  assign core_rc_tuser_sop0_lower = core_rc_tuser_reg_lower_user_clk_int[32];
  assign core_rc_tuser_sop1_lower = core_rc_tuser_reg_lower_user_clk_int[33];
  assign core_rc_tuser_eop0_lower = core_rc_tuser_reg_lower_user_clk_int[34];
  assign core_rc_tuser_eop1_lower = core_rc_tuser_reg_lower_user_clk_int[38];

  assign core_rc_tuser_sop0_upper = core_rc_tuser_reg_upper_user_clk_int[32];
  assign core_rc_tuser_sop1_upper = core_rc_tuser_reg_upper_user_clk_int[33];
  assign core_rc_tuser_eop0_upper = core_rc_tuser_reg_upper_user_clk_int[34];
  assign core_rc_tuser_eop1_upper = core_rc_tuser_reg_upper_user_clk_int[38];

  always @(posedge user_clk_i)
    if (~reset_n_user_clk_i)
      core_rc_pkt_in_progress <= #TCQ 1'b0;
    else if (link_down_reset_i)
      core_rc_pkt_in_progress <= #TCQ 1'b0;
    else
      if (~core_rc_pkt_in_progress)
    begin
      case({core_rc_tvalid_reg_upper_user_clk, core_rc_tvalid_reg_lower_user_clk})
        2'b00:
          begin
          end
        2'b01:
          begin
        core_rc_pkt_in_progress <= #TCQ 1'b0;
          end
        2'b10:
          begin
        core_rc_pkt_in_progress <= #TCQ ~core_rc_tuser_eop0_upper |
                       (core_rc_tuser_sop1_upper & ~core_rc_tuser_eop1_upper);
          end
        2'b11:
          begin
        core_rc_pkt_in_progress <= #TCQ ((~core_rc_tuser_eop0_lower |
                          (core_rc_tuser_sop1_lower & ~core_rc_tuser_eop1_lower)) &
                          (~core_rc_tuser_eop0_upper |
                           (core_rc_tuser_sop0_upper & ~core_rc_tuser_eop1_upper))) |
                       (((core_rc_tuser_eop0_lower & ~core_rc_tuser_sop1_lower) |
                         core_rc_tuser_eop1_lower) &
                        (~core_rc_tuser_eop0_upper |
                         (core_rc_tuser_sop1_upper & ~core_rc_tuser_eop1_upper)));
          end // case: 2'b11
      endcase // case({core_rc_tvalid_reg_upper_user_clk, core_rc_tvalid_reg_lower_user_clk})
    end // if (~core_rc_pkt_in_progress)
      else
      begin      
      case({core_rc_tvalid_reg_upper_user_clk, core_rc_tvalid_reg_lower_user_clk})
        2'b00:
          begin
          end
        2'b01:
          begin
        core_rc_pkt_in_progress <= #TCQ 1'b0;
          end
        2'b10:
          begin
        // Invalid case
        core_rc_pkt_in_progress <= #TCQ 1'b0;
          end
         2'b11:
           begin
         core_rc_pkt_in_progress <= #TCQ ((~core_rc_tuser_eop0_lower |
                           (core_rc_tuser_sop0_lower & ~core_rc_tuser_eop1_lower)) &
                          (~core_rc_tuser_eop0_upper |
                           (core_rc_tuser_sop0_upper & ~core_rc_tuser_eop1_upper))) |
                        (((core_rc_tuser_eop0_lower & ~core_rc_tuser_sop0_lower) |
                          core_rc_tuser_eop1_lower) &
                         (~core_rc_tuser_eop0_upper |
                          (core_rc_tuser_sop1_upper & ~core_rc_tuser_eop1_upper)));
           end // case: 2'b11
      endcase // case({core_rc_tvalid_reg_upper_user_clk, core_rc_tvalid_reg_lower_user_clk})
    end // else: !if(~core_rc_pkt_in_progress)

  assign core_rc_pkt_in_progress_upper = ~core_rc_tvalid_reg_lower_user_clk? 1'b0:
                     core_rc_pkt_in_progress? (~core_rc_tuser_eop0_lower |
                                   (core_rc_tuser_sop0_lower & ~core_rc_tuser_eop1_lower)):
                     (~core_rc_tuser_eop0_lower |
                      (core_rc_tuser_sop1_lower & ~core_rc_tuser_eop1_lower));

  assign core_rc_tuser_reg_sop0_ptr_lower = ~attr_straddle_en_i? 1'b0:
     core_rc_pkt_in_progress? 
     core_rc_tvalid_reg_lower_user_clk & core_rc_tuser_sop0_lower : 1'b0;

  assign core_rc_tuser_reg_sop0_ptr_upper = ~attr_straddle_en_i? 1'b0:
     core_rc_pkt_in_progress_upper? 
         core_rc_tvalid_reg_upper_user_clk & core_rc_tuser_sop0_upper : 1'b0;
  
   // Write data into FIFO using 250 MHz user_clk

  generate
    if (PARITY_ENABLE)
      assign fifo_in_data =
          {
       core_rc_tvalid_reg_upper_user_clk,
       core_rc_tlast_reg_upper_user_clk,
       core_rc_tuser_reg_sop0_ptr_upper, 
       core_rc_tuser_reg_upper_user_clk_int,
       core_rc_tkeep_reg_upper_user_clk,
       core_rc_tdata_reg_upper_user_clk,
       core_rc_tvalid_reg_lower_user_clk,
       core_rc_tlast_reg_lower_user_clk,
       core_rc_tuser_reg_sop0_ptr_lower, 
       core_rc_tuser_reg_lower_user_clk_int,
       core_rc_tkeep_reg_lower_user_clk,
       core_rc_tdata_reg_lower_user_clk
       };
    else
      assign fifo_in_data =
          {
       core_rc_tvalid_reg_upper_user_clk,
       core_rc_tlast_reg_upper_user_clk,
       core_rc_tuser_reg_sop0_ptr_upper, 
       core_rc_tuser_reg_upper_user_clk_int[42:0],
       core_rc_tkeep_reg_upper_user_clk,
       core_rc_tdata_reg_upper_user_clk,
       core_rc_tvalid_reg_lower_user_clk,
       core_rc_tlast_reg_lower_user_clk,
       core_rc_tuser_reg_sop0_ptr_lower, 
       core_rc_tuser_reg_lower_user_clk_int[42:0],
       core_rc_tkeep_reg_lower_user_clk,
       core_rc_tdata_reg_lower_user_clk
       };
  endgenerate

   // Generate ready to core in the user_clk2 domain
   always @(posedge user_clk2_i)
     if (~reset_n_user_clk2_i)
       begin
      core_rc_tready_user_clk2 <= #TCQ 1'b0;
      core_rc_tready_reg <= #TCQ {AXI4_CORE_RC_TREADY_WIDTH{1'b0}};
       end
     else
       begin
             core_rc_tready_user_clk2 <= #TCQ ~fifo_almost_full_user_clk;
      core_rc_tready_reg <= #TCQ {AXI4_CORE_RC_TREADY_WIDTH{~fifo_almost_full_user_clk}};
       end

   assign core_rc_tready_o = core_rc_tready_reg;
 

   // Main FIFO instance
   xp4_usp_smsw_512b_sync_fifo #
     (
      .TCQ(TCQ),
      .IMPL_TARGET(IMPL_TARGET),
      .AXISTEN_IF_EXT_512_INTFC_RAM_STYLE(AXISTEN_IF_EXT_512_INTFC_RAM_STYLE),
      .FIFO_WIDTH(FIFO_WIDTH),
      .FIFO_DEPTH(8),
      .FIFO_ALMOST_FULL_THRESHOLD(5)
      )
     pcie_4_0_512b_sync_fifo_blk
       (
        .clk_i(user_clk_i),
        .reset_n_i(reset_n_user_clk_i),
        .link_down_reset_i(link_down_reset_i),
    .write_data_i(fifo_in_data),
    .write_en_i(fifo_in_data_valid),
    .read_en_i(fifo_read_en),
    .read_data_o(fifo_read_data),
    .read_data_valid_o(fifo_read_data_valid),
    .fifo_almost_full(fifo_almost_full_user_clk)
    );
   
   // Read-side logic

   assign read_sop0_lower = fifo_read_data[TUSER_LOWER_OFFSET + 32];
   assign read_sop1_lower = fifo_read_data[TUSER_LOWER_OFFSET + 33];
   assign  read_eop0_lower = fifo_read_data[TUSER_LOWER_OFFSET + 34];
   assign  read_eop1_lower = fifo_read_data[TUSER_LOWER_OFFSET + 38];
   assign read_discontinue_lower = fifo_read_data[TUSER_LOWER_OFFSET + 42];

   assign read_sop0_upper = fifo_read_data[TUSER_UPPER_OFFSET + 32];
   assign read_sop1_upper = fifo_read_data[TUSER_UPPER_OFFSET + 33];
   assign  read_eop0_upper = fifo_read_data[TUSER_UPPER_OFFSET + 34];
   assign  read_eop1_upper = fifo_read_data[TUSER_UPPER_OFFSET + 38];
   assign read_discontinue_upper = fifo_read_data[TUSER_UPPER_OFFSET + 42];

  generate
    if (PARITY_ENABLE)
      begin
    assign read_sop0_ptr_lower = fifo_read_data[TUSER_LOWER_OFFSET + AXI4_CORE_RC_TUSER_WIDTH];
    assign read_sop0_ptr_upper = fifo_read_data[TUSER_UPPER_OFFSET + AXI4_CORE_RC_TUSER_WIDTH];
    assign read_tlast_lower = fifo_read_data[AXI4_CORE_DATA_WIDTH + AXI4_CORE_RC_TKEEP_WIDTH +
                         AXI4_CORE_RC_TUSER_WIDTH+1];
    assign read_tlast_upper = fifo_read_data[AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_RC_TKEEP_WIDTH*2 +
                         (AXI4_CORE_RC_TUSER_WIDTH+1)*2 +2];
      end
    else
      begin
    assign read_sop0_ptr_lower = fifo_read_data[TUSER_LOWER_OFFSET + AXI4_CORE_RC_TUSER_WIDTH-32];
    assign read_sop0_ptr_upper = fifo_read_data[TUSER_UPPER_OFFSET + AXI4_CORE_RC_TUSER_WIDTH-64];
    assign read_tlast_lower = fifo_read_data[AXI4_CORE_DATA_WIDTH + AXI4_CORE_RC_TKEEP_WIDTH +
                         (AXI4_CORE_RC_TUSER_WIDTH+1) -32];
    assign read_tlast_upper = fifo_read_data[AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_RC_TKEEP_WIDTH*2 +
                         (AXI4_CORE_RC_TUSER_WIDTH+1)*2 +2 -64];
      end // else: !if(PARITY_ENABLE)
  endgenerate

    assign        read_data_valid_lower = fifo_read_data[FIFO_WIDTH/2-1] & fifo_read_data_valid;
    assign        read_data_valid_upper = fifo_read_data[FIFO_WIDTH-1] & fifo_read_data_valid;

  assign        read_sop_upper = read_sop0_upper;

  assign        read_eop_lower = ~attr_straddle_en_i? read_tlast_lower:
           ~read_sop0_lower? // No new TLP starting
           read_eop0_lower:
           (read_sop0_lower & ~read_sop0_ptr_lower)? // New TLP starting on DW 0
           ((read_eop0_lower & ~read_sop1_lower) | read_eop1_lower):
           (read_sop0_lower & read_sop0_ptr_lower)? // TLP contiuning from last beat, new TLP starting on DW 4
           read_eop1_lower: 1'b0;
  
  assign        read_eop_upper = ~attr_straddle_en_i? read_tlast_upper:
           ~read_sop0_upper? // No new TLP starting
           read_eop0_upper:
           (read_sop0_upper & ~read_sop0_ptr_upper)? // New TLP starting on DW 0
           ((read_eop0_upper & ~read_sop1_upper) | read_eop1_upper):
           (read_sop0_upper & read_sop0_ptr_upper)? // TLP contiuning from last beat, new TLP starting on DW 4
           read_eop1_upper: 1'b0;

   // Read State Machine States
   //
   // IDLE: Currently not forwarding a packet.  Read data register is either empty, or contains the last beat of a packet.
   // EXPECT_NEW_WORD: Currently forwarding a packet, and there is no data saved from a previous beat
   // SEND_SAVED_HALF_WORD: There is a half-word saved from a previous beat in the saved data register.
   // WAIT_FOR_UPPER_HALF: There is a half-word saved from a previous beat in the read data register which does not end with an EOP.
   
   always @(posedge user_clk_i)
     if (~reset_n_user_clk_i)
       begin
      read_data_valid_reg <= #TCQ 2'b00;
      read_state <= #TCQ IDLE;
       end
     else if (link_down_reset_i)
       begin
      read_data_valid_reg <= #TCQ 2'b00;
      read_state <= #TCQ IDLE;
       end
     else
    case(read_state)
      IDLE:
        begin
           // IDLE: Currently not forwarding a packet.  Read data register is either empty, or contains the last beat of a packet.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if (read_data_valid_lower)
              // New TLP starting in the lower half of the incoming word.
              // Update the lower half of the data register with the lower half of the incoming word.
              begin
             if (read_data_valid_upper)
               // Both halves of the incoming word have valid data in them.
               begin
                  // If straddle is not enabled and the packet in the upper half is a new one,
                  // Save it for next cycle.
                  // Also, if the packet in the lower half ends with an error, do not fill the upper half.
                  if ((~attr_straddle_en_i & read_sop_upper)|
                  read_discontinue_lower)
                begin
                   read_data_valid_reg <= #TCQ 2'b01;
                   read_state <= #TCQ SEND_SAVED_HALF_WORD;
                end
                  else
                begin
                   read_data_valid_reg <= #TCQ 2'b11;
                  if (read_eop_upper)
                     read_state <= #TCQ IDLE;
                   else
                     read_state <= #TCQ EXPECT_NEW_WORD;
                end // else: !if(~attr_straddle_en_i & read_sop_upper)
               end // if (read_data_valid_upper)
             else
               begin
                  // New TLP started in the lower half, but there is no valid data in the upper half.
                  if (read_eop_lower)
                // We have a complete TLP in the lower half, send it.
                begin
                   read_data_valid_reg <= #TCQ 2'b01;
                   read_state <= #TCQ IDLE;
                end
                  else
                begin
                   // Wait for more data to fill upper half of read data register.
                   read_data_valid_reg <= #TCQ 2'b00;
                   read_state <= #TCQ WAIT_FOR_UPPER_HALF;
                end // else: !if(read_eop_lower)
               end // else: !if(read_data_valid_upper)
              end // if (read_data_valid_lower)
            else
              if (read_data_valid_upper)
            begin
               // No valid data in the lower half of the incoming word, but there is a packet starting in the upper half.
               if (read_eop_upper)
                 // We have a complete packet, send it in the lower half.
                 begin
                read_data_valid_reg <= #TCQ 2'b01;
                read_state <= #TCQ IDLE;
                 end
               else
                 begin
                // Save the upper half of the incoming word
                // and wait for more data.
                read_data_valid_reg <= #TCQ 2'b00;
                read_state <= #TCQ WAIT_FOR_UPPER_HALF;
                 end // else: !if(read_eop_upper)
            end // if (read_data_valid_upper)
              else
            // No valid data from FIFO
            begin
               if (output_mux_ready)
                 read_data_valid_reg <= #TCQ 2'b00;
               read_state <= #TCQ IDLE;
            end // else: !if(read_data_valid_upper)
         end // if ((read_data_valid_reg == 2'b00) | output_mux_ready)
        end // case: IDLE
      
      EXPECT_NEW_WORD:
        begin
           // Currently forwarding a packet.  There is no saved data.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if (read_data_valid_lower)
              // New data starting in the lower half of the incoming word.
              // Update the lower half of the data register with the lower half of the incoming word.
              begin
             if (read_data_valid_upper)
               // Both halves of the incoming word have valid data in them.
               begin
                  // If straddle is not enabled and the packet in the upper half is a new one,
                  // Save it for next cycle.
                  // Also, if the packet in the lower half ends with an error, do not fill the upper half.
                  if ((~attr_straddle_en_i & read_sop_upper)|
                  read_discontinue_lower)
                begin
                   read_data_valid_reg <= #TCQ 2'b01;
                   read_state <= #TCQ SEND_SAVED_HALF_WORD;
                end
                  else
                begin
                   read_data_valid_reg <= #TCQ 2'b11;
                  if (read_eop_upper)
                     read_state <= #TCQ IDLE;
                  else
                     read_state <= #TCQ EXPECT_NEW_WORD;
                end // else: !if((~attr_straddle_en_i & read_sop_upper)|...
               end // if (read_data_valid_upper)
             else
               begin
                  // Valid data in the lower half, but no valid data in the upper half.
                  if (read_eop_lower)
                // We have the packet ending in the lower half, send it.
                begin
                   read_data_valid_reg <= #TCQ 2'b01;
                   read_state <= #TCQ IDLE;
                end
                  else
                begin
                   // Wait for more data to fill upper half of read data register.
                   read_data_valid_reg <= #TCQ 2'b00;
                   read_state <= #TCQ WAIT_FOR_UPPER_HALF;
                end // else: !if(read_eop_lower)
               end // else: !if(read_data_valid_upper)
              end // if (read_data_valid_lower)
            else
              if (read_data_valid_upper)
            begin
               // No valid data in the lower half of the incoming word, but there is data in the upper half.
               if (read_eop_upper)
                 // We have a complete packet, send it in the lower half.
                 begin
                read_data_valid_reg <= #TCQ 2'b01;
                read_state <= #TCQ IDLE;
                 end
               else
                 begin
                // Save the upper half of the incoming word
                // and wait for more data.
                read_data_valid_reg <= #TCQ 2'b00;
                read_state <= #TCQ WAIT_FOR_UPPER_HALF;
                 end // else: !if(read_eop_upper)
            end // if (read_data_valid_upper)
              else
            // No valid data from FIFO
            begin
               if (output_mux_ready)
                 read_data_valid_reg <= #TCQ 2'b00;
               read_state <= #TCQ EXPECT_NEW_WORD;
            end // else: !if(read_data_valid_upper)
         end // if ((read_data_valid_reg == 2'b00) | output_mux_ready)
        end // case: EXPECT_NEW_WORD

      SEND_SAVED_HALF_WORD:
        begin
           // There is a half-word saved from a previous beat in the saved data register.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if ((~attr_straddle_en_i & saved_eop) | saved_err)
              // Saved data is the last beat of a packet and straddle is disabled.
              // Do not fill the upper half of read data register.
              begin
            read_data_valid_reg <= #TCQ 2'b01;
            read_state <= #TCQ IDLE;
              end
            else
              if (read_data_valid_lower)
            // New data starting in the lower half of the incoming word.
            // Update the upper half of the data register with the lower half of the incoming word.
            begin
               if (read_data_valid_upper)
                 // Both halves of the incoming word have valid data in them.
                 begin
                read_data_valid_reg <= #TCQ 2'b11;
                read_state <= #TCQ SEND_SAVED_HALF_WORD;
                 end
               else
                 begin
                read_data_valid_reg <= #TCQ 2'b11;
                if (read_eop_lower)
                  read_state <= #TCQ IDLE;
                else
                  read_state <= #TCQ EXPECT_NEW_WORD;
                 end // else: !if(read_data_valid_upper)
            end // if (read_data_valid_lower)
              else
            if (read_data_valid_upper)
              begin
                 // No valid data in the lower half of the incoming word, but there is data in the upper half.
                 if (read_eop_upper)
                   // We have a complete packet, send it in the upper half.
                   begin
                  read_data_valid_reg <= #TCQ 2'b11;
                  read_state <= #TCQ IDLE;
                   end
                 else
                   begin
                  read_data_valid_reg <= #TCQ 2'b11;
                  read_state <= #TCQ EXPECT_NEW_WORD;
                   end // else: !if(read_eop_upper)
              end // if (read_data_valid_upper)
            else
              // No valid data from FIFO
              begin
                read_data_valid_reg <= #TCQ 2'b01;
                read_state <= #TCQ IDLE;
              end // else: !if(read_data_valid_upper)
         end // if ((read_data_valid_reg == 2'b00) | output_mux_ready)
        end // case: SEND_SAVED_HALF_WORD

      WAIT_FOR_UPPER_HALF:
        begin
           // There is a half-word saved from a previous beat in the read data register which does not end with an EOP.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if (read_data_valid_lower)
              // New data starting in the lower half of the incoming word.
              // Update the upper half of the data register with the lower half of the incoming word.
              begin
             read_data_valid_reg <= #TCQ 2'b11;
             if (read_data_valid_upper)
               // Both halves of the incoming word have valid data in them.
               begin
                 if (read_eop_upper)
                   read_state <= #TCQ SEND_SAVED_HALF_WORD;
                 else
                   read_state <= #TCQ WAIT_FOR_UPPER_HALF;
               end
             else
               begin
                 if (read_eop_lower)
                   read_state <= #TCQ IDLE;
                 else
                   read_state <= #TCQ EXPECT_NEW_WORD;
               end // else: !if(read_data_valid_upper)
              end // if (read_data_valid_lower)
            else
              if (read_data_valid_upper)
            begin
               // No valid data in the lower half of the incoming word, but there is data in the upper half.
               read_data_valid_reg <= #TCQ 2'b11;
               if (read_eop_upper)
                 read_state <= #TCQ IDLE;
               else
                 read_state <= #TCQ EXPECT_NEW_WORD;
            end // if (read_data_valid_upper)
              else
            begin
               read_data_valid_reg <= #TCQ 2'b00;
               read_state <= #TCQ WAIT_FOR_UPPER_HALF;
            end // else: !if(read_data_valid_upper)
         end // if ((read_data_valid_reg == 2'b00) | output_mux_ready)
        end // case: WAIT_FOR_UPPER_HALF
    endcase // case(read_state)

   always @(posedge user_clk_i)
     if (~reset_n_user_clk_i)
       begin
      read_data_reg <= #TCQ {FIFO_WIDTH{1'b0}};
      saved_data_reg <= #TCQ {FIFO_WIDTH/2{1'b0}};
      saved_eop <= #TCQ 1'b0;
      saved_err <= #TCQ 1'b0;
       end
     else
    case(read_state)
      IDLE:
        begin
           // IDLE: Currently not forwarding a packet.  Read data register is either empty, or contains the last beat of a packet.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if (read_data_valid_lower)
              read_data_reg[FIFO_WIDTH/2-1:0] <= #TCQ fifo_read_data[FIFO_WIDTH/2-1:0];
            else
              read_data_reg[FIFO_WIDTH/2-1:0] <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
            read_data_reg[FIFO_WIDTH-1: FIFO_WIDTH/2] <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
            saved_data_reg <= #TCQ fifo_read_data[FIFO_WIDTH-1:FIFO_WIDTH/2];
            saved_eop <= #TCQ read_eop_upper;
            saved_err <= #TCQ read_discontinue_upper;
         end
        end // case: IDLE

      EXPECT_NEW_WORD:
        begin
           // Currently not forwarding a packet.  
           // Read data register is either empty, or contains the last beat of a packet.           
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if (read_data_valid_lower)
              read_data_reg[FIFO_WIDTH/2-1:0] <= #TCQ fifo_read_data[FIFO_WIDTH/2-1:0];
            else
              read_data_reg[FIFO_WIDTH/2-1:0] <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
            read_data_reg[FIFO_WIDTH-1: FIFO_WIDTH/2] <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
            saved_data_reg <= #TCQ fifo_read_data[FIFO_WIDTH-1:FIFO_WIDTH/2];
            saved_eop <= #TCQ read_eop_upper;
            saved_err <= #TCQ read_discontinue_upper;
         end
        end // case: EXPECT_NEW_WORD
      
      SEND_SAVED_HALF_WORD:
        begin
           // There is a half-word saved from a previous beat in the saved data register.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            read_data_reg[FIFO_WIDTH/2-1:0] <= #TCQ saved_data_reg[FIFO_WIDTH/2-1: 0];
            if (read_data_valid_lower)
              read_data_reg[FIFO_WIDTH-1: FIFO_WIDTH/2] <= #TCQ fifo_read_data[FIFO_WIDTH/2-1: 0];
            else
              read_data_reg[FIFO_WIDTH-1: FIFO_WIDTH/2] <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
            

            if ((~attr_straddle_en_i & saved_eop) | saved_err)
              // Save incoming data for next cycle.
              begin
             if (read_data_valid_lower)
               begin
                  saved_data_reg <= #TCQ fifo_read_data[FIFO_WIDTH/2-1: 0];
                  saved_eop <= #TCQ read_eop_lower;
                  saved_err <= #TCQ read_discontinue_lower;
               end
             else
               begin
                  saved_data_reg <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
                  saved_eop <= #TCQ read_eop_upper;
                  saved_err <= #TCQ read_discontinue_upper;
               end
              end
            else
              begin
             saved_data_reg <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
             saved_eop <= #TCQ read_eop_upper;
             saved_err <= #TCQ read_discontinue_upper;
              end // else: !if((~attr_straddle_en_i & saved_eop) | saved_err)
         end // if ((read_data_valid_reg == 2'b00) | output_mux_ready)
        end // case: SEND_SAVED_HALF_WORD
      WAIT_FOR_UPPER_HALF:
        begin
           // There is a half-word saved from a previous beat in the read data register which does not end with an EOP.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
           read_data_reg[FIFO_WIDTH/2-1:0] <= #TCQ saved_data_reg[FIFO_WIDTH/2-1:0];
            if (read_data_valid_lower)
              read_data_reg[FIFO_WIDTH-1: FIFO_WIDTH/2] <= #TCQ fifo_read_data[FIFO_WIDTH/2-1: 0];
            else
              read_data_reg[FIFO_WIDTH-1: FIFO_WIDTH/2] <= #TCQ {FIFO_WIDTH/2{1'b0}};
              // Save incoming data for next cycle.
            saved_data_reg <= #TCQ fifo_read_data[FIFO_WIDTH-1: FIFO_WIDTH/2];
            saved_eop <= #TCQ read_eop_upper;
            saved_err <= #TCQ read_discontinue_upper;
         end
        end // case: WAIT_FOR_UPPER_HALF
    endcase // case(read_state)
         
   // Generate upstream ready
   always @(*)
     begin
    case(read_state)
      IDLE:
        begin
           fifo_read_en = (read_data_valid_reg == 2'b00) | output_mux_ready;
        end
      
      EXPECT_NEW_WORD:
        begin
           fifo_read_en = (read_data_valid_reg == 2'b00) | output_mux_ready;
        end

      SEND_SAVED_HALF_WORD:
        begin
           // There is a half-word saved from a previous beat in the saved data register.
           if ((read_data_valid_reg == 2'b00) | output_mux_ready)
         begin
            if ((~attr_straddle_en_i & saved_eop) | saved_err)
              // Saved data is the last beat of a packet and straddle is disabled.
              // Do not fill the upper half of read data register.
              fifo_read_en = 1'b0;
            else
              fifo_read_en = 1'b1;
         end
           else
         fifo_read_en = 1'b0;
        end // case: SEND_SAVED_HALF_WORD

      WAIT_FOR_UPPER_HALF:
        begin
           // There is a half-word saved from a previous beat in the read data register which does not end with an EOP.
           fifo_read_en = (read_data_valid_reg == 2'b00) | output_mux_ready;
        end
    endcase // case(read_state)
     end // always @ (*)
   
   assign read_data_reg_byte_en_lower = read_data_reg[TUSER_LOWER_OFFSET +31:
                                 TUSER_LOWER_OFFSET];
   assign read_data_reg_sop0_lower = read_data_reg[TUSER_LOWER_OFFSET + 32];
  assign  read_data_reg_sop1_lower = attr_straddle_en_i? read_data_reg[TUSER_LOWER_OFFSET + 33]: 1'b0;
   assign read_data_reg_eop0_lower = attr_straddle_en_i? read_data_reg[TUSER_LOWER_OFFSET + 34]:
      read_data_reg_tlast_lower;
   assign read_data_reg_eop0_ptr_lower[2:0] = read_data_reg[TUSER_LOWER_OFFSET + 37:
                                TUSER_LOWER_OFFSET + 35];
  assign  read_data_reg_eop1_lower = attr_straddle_en_i? read_data_reg[TUSER_LOWER_OFFSET + 38]: 1'b0;
   assign read_data_reg_eop1_ptr_lower[2:0] = attr_straddle_en_i? read_data_reg[TUSER_LOWER_OFFSET + 41:
                                        TUSER_LOWER_OFFSET + 39]: 3'd0;
   assign read_data_reg_discontinue_lower = read_data_reg[TUSER_LOWER_OFFSET + 42];

  generate
    if (PARITY_ENABLE)
      begin
    assign read_data_reg_parity_lower = read_data_reg[TUSER_LOWER_OFFSET + 74:   
                                   TUSER_LOWER_OFFSET + 43];
    assign read_data_reg_sop0_ptr_lower = read_data_reg[TUSER_LOWER_OFFSET + 75];
      end
    else
      begin
    assign read_data_reg_parity_lower = 32'd0;
    assign read_data_reg_sop0_ptr_lower = read_data_reg[TUSER_LOWER_OFFSET + 43];
      end // else: !if(PARITY_ENABLE)
  endgenerate
  
  assign     read_data_reg_byte_en_upper = read_data_reg[TUSER_UPPER_OFFSET +31:
                                 TUSER_UPPER_OFFSET];
   assign read_data_reg_sop0_upper = read_data_reg[TUSER_UPPER_OFFSET + 32];
  assign  read_data_reg_sop1_upper = attr_straddle_en_i? read_data_reg[TUSER_UPPER_OFFSET + 33]: 1'b0;
   assign read_data_reg_eop0_upper = attr_straddle_en_i? read_data_reg[TUSER_UPPER_OFFSET + 34]:
      read_data_reg_tlast_upper;
   assign read_data_reg_eop0_ptr_upper[2:0] = read_data_reg[TUSER_UPPER_OFFSET + 37:
                                TUSER_UPPER_OFFSET + 35];
   assign read_data_reg_eop1_upper = attr_straddle_en_i? read_data_reg[TUSER_UPPER_OFFSET + 38]: 1'b0;
   assign read_data_reg_eop1_ptr_upper[2:0] = attr_straddle_en_i? read_data_reg[TUSER_UPPER_OFFSET + 41:
                                        TUSER_UPPER_OFFSET + 39]: 3'd0;
   assign read_data_reg_discontinue_upper = read_data_reg[TUSER_UPPER_OFFSET + 42];

  generate
    if (PARITY_ENABLE)
      begin
    assign read_data_reg_parity_upper = read_data_reg[TUSER_UPPER_OFFSET + 74:   
                                   TUSER_UPPER_OFFSET + 43];
    assign read_data_reg_sop0_ptr_upper = read_data_reg[TUSER_UPPER_OFFSET + 75];
      end
    else
      begin
    assign read_data_reg_parity_upper = 32'd0;
    assign read_data_reg_sop0_ptr_upper = read_data_reg[TUSER_UPPER_OFFSET + 43];
      end // else: !if(PARITY_ENABLE)
  endgenerate

  generate
    if (PARITY_ENABLE)
      begin
    assign  read_data_reg_tlast_lower = read_data_reg[AXI4_CORE_DATA_WIDTH + AXI4_CORE_RC_TKEEP_WIDTH +
                              AXI4_CORE_RC_TUSER_WIDTH+1];
    assign     read_data_reg_tlast_upper = read_data_reg[AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_RC_TKEEP_WIDTH*2 +
                              (AXI4_CORE_RC_TUSER_WIDTH+1)*2 +2];
      end
    else
      begin
    assign  read_data_reg_tlast_lower = read_data_reg[AXI4_CORE_DATA_WIDTH + AXI4_CORE_RC_TKEEP_WIDTH +
                              AXI4_CORE_RC_TUSER_WIDTH+1 -32];
    assign     read_data_reg_tlast_upper = read_data_reg[AXI4_CORE_DATA_WIDTH*2 + AXI4_CORE_RC_TKEEP_WIDTH*2 +
                              (AXI4_CORE_RC_TUSER_WIDTH+1)*2 +2 -64];
      end // else: !if(PARITY_ENABLE)
  endgenerate

   assign read_data_out_byte_en[31:0] = read_data_valid_reg[0]? read_data_reg_byte_en_lower: 32'd0;
   assign read_data_out_byte_en[63:32] = read_data_valid_reg[1]? read_data_reg_byte_en_upper: 32'd0;

  assign  read_data_out_is_sop[0] = ((read_data_valid_reg[0] & (read_data_reg_sop0_lower | 
                                read_data_reg_sop1_lower))) |
      ((read_data_valid_reg[1] & (read_data_reg_sop0_upper | read_data_reg_sop1_upper)));
  
  assign  read_data_out_is_sop[1] = (read_data_valid_reg[0] & read_data_reg_sop1_lower) | 
      (read_data_valid_reg[1] & read_data_reg_sop1_upper) | 
      (read_data_valid_reg[0] & read_data_reg_sop0_lower & read_data_valid_reg[1] &
       read_data_reg_sop0_upper);

  assign  read_data_out_is_sop[2] = read_data_valid_reg[0] & read_data_valid_reg[1] & 
      ((read_data_reg_sop1_lower & read_data_reg_sop0_upper) |
       (read_data_reg_sop0_lower & read_data_reg_sop1_upper));
  
  assign  read_data_out_is_sop[3] = read_data_valid_reg[0] & read_data_valid_reg[1] & 
      read_data_reg_sop1_lower & read_data_reg_sop1_upper;

  assign  read_data_out_is_sop0_ptr[1:0] = (read_data_valid_reg[0] & read_data_reg_sop0_lower)?
      {1'b0, read_data_reg_sop0_ptr_lower}:
      (read_data_valid_reg[0] & read_data_reg_sop1_lower)? 2'd1:
      (read_data_valid_reg[1] & read_data_reg_sop0_upper)?
      {1'b1, read_data_reg_sop0_ptr_upper}:
      (read_data_valid_reg[1] & read_data_reg_sop1_upper)? 2'd3: 2'd0;
  assign  read_data_out_is_sop1_ptr[1:0] = (read_data_valid_reg[0] & read_data_reg_sop1_lower)? 4'd1:
      (read_data_valid_reg[0] & read_data_valid_reg[1] & read_data_reg_sop0_lower &
       read_data_reg_sop0_upper)? {1'b1, read_data_reg_sop0_ptr_upper}:
      (read_data_valid_reg[1] & read_data_reg_sop0_upper &
       read_data_reg_sop1_upper)? 2'd3: 2'd0;
    assign  read_data_out_is_sop2_ptr[1:0] = (read_data_valid_reg[0] & read_data_valid_reg[1] & 
                          read_data_reg_sop1_lower & read_data_reg_sop0_upper)? 
        {1'b1, read_data_reg_sop0_ptr_upper}:
        (read_data_valid_reg[0] & read_data_valid_reg[1] & 
         read_data_reg_sop0_lower & read_data_reg_sop1_upper)? 2'd3: 2'd0;
  assign    read_data_out_is_sop3_ptr[1:0] = (read_data_valid_reg[0] & read_data_valid_reg[1] & 
                          read_data_reg_sop1_lower & read_data_reg_sop1_upper)? 2'd3: 2'd0;

  assign  read_data_out_is_eop[0] = ((read_data_valid_reg[0] & (read_data_reg_eop0_lower | 
                                read_data_reg_eop1_lower))) |
      ((read_data_valid_reg[1] & (read_data_reg_eop0_upper | read_data_reg_eop1_upper)));

  assign  read_data_out_is_eop0_ptr[3:0] = (read_data_valid_reg[0] & read_data_reg_eop0_lower)?
       {1'b0, read_data_reg_eop0_ptr_lower[2:0]}:
      (read_data_valid_reg[0] & read_data_reg_eop1_lower)?
       {1'b0, read_data_reg_eop1_ptr_lower[2:0]}:
      (read_data_valid_reg[1] & read_data_reg_eop0_upper)?
       {1'b1, read_data_reg_eop0_ptr_upper[2:0]}:
      (read_data_valid_reg[1] & read_data_reg_eop1_upper)?
       {1'b1, read_data_reg_eop1_ptr_upper[2:0]}: 4'd0;
  
  assign  read_data_out_is_eop[1] = (read_data_valid_reg[0] & read_data_reg_eop1_lower) | 
      (read_data_valid_reg[1] & read_data_reg_eop1_upper) | 
      (read_data_valid_reg[0] & read_data_reg_eop0_lower & read_data_valid_reg[1] &
       read_data_reg_eop0_upper);
  assign  read_data_out_is_eop1_ptr[3:0] = (read_data_valid_reg[0] & read_data_reg_eop1_lower)?
       {1'b0, read_data_reg_eop1_ptr_lower[2:0]}:
      (read_data_valid_reg[0] & read_data_reg_eop0_lower & 
       read_data_valid_reg[1] & read_data_reg_eop0_upper)?
       {1'b1, read_data_reg_eop0_ptr_upper[2:0]}:
      (read_data_valid_reg[1] & read_data_reg_eop1_upper)?
      {1'b1, read_data_reg_eop1_ptr_upper[2:0]}: 4'd0;

  assign  read_data_out_is_eop[2] = read_data_valid_reg[0] & read_data_valid_reg[1] & 
      ((read_data_reg_eop1_lower & read_data_reg_eop0_upper) |
       (read_data_reg_eop0_lower & read_data_reg_eop1_upper));
  assign  read_data_out_is_eop2_ptr[3:0] = (read_data_valid_reg[0] & read_data_valid_reg[1] & 
                        read_data_reg_eop1_lower & read_data_reg_eop0_upper)?
       {1'b1, read_data_reg_eop0_ptr_upper[2:0]}:
      (read_data_valid_reg[0] & read_data_valid_reg[1] & 
       read_data_reg_eop0_lower & read_data_reg_eop1_upper)?
       {1'b1, read_data_reg_eop1_ptr_upper[2:0]}: 4'd0;
  assign  read_data_out_is_eop[3] = read_data_valid_reg[0] & read_data_valid_reg[1] & 
      read_data_reg_eop1_lower & read_data_reg_eop1_upper;
  assign  read_data_out_is_eop3_ptr[3:0] = (read_data_valid_reg[0] & read_data_valid_reg[1] & 
                        read_data_reg_eop1_lower & read_data_reg_eop1_upper)?
      {1'b1, read_data_reg_eop1_ptr_upper[2:0]}: 4'd0;

   assign read_data_out_discontinue = (read_data_valid_reg[0] & read_data_reg_discontinue_lower) |
      (read_data_valid_reg[1] & read_data_reg_discontinue_upper);      

   assign read_data_out_parity[31:0] = read_data_valid_reg[0]? read_data_reg_parity_lower: 32'd0;
   assign read_data_out_parity[63:32] = read_data_valid_reg[1]? read_data_reg_parity_upper: 32'd0;  

   assign read_data_out_tuser = {
                 read_data_out_parity[63:0],
                 read_data_out_discontinue,
                 read_data_out_is_eop3_ptr[3:0],
                 read_data_out_is_eop2_ptr[3:0],
                 read_data_out_is_eop1_ptr[3:0],
                 read_data_out_is_eop0_ptr[3:0],
                 read_data_out_is_eop[3:0],
                 read_data_out_is_sop3_ptr[1:0],
                 read_data_out_is_sop2_ptr[1:0],
                 read_data_out_is_sop1_ptr[1:0],
                 read_data_out_is_sop0_ptr[1:0],
                 read_data_out_is_sop[3:0],
                 read_data_out_byte_en[63:0]
                 };

   assign read_data_out_tdata[AXI4_USER_DATA_WIDTH/2-1:0] = read_data_valid_reg[0]? read_data_reg[AXI4_CORE_DATA_WIDTH-1:0]:
      {AXI4_USER_DATA_WIDTH/2{1'b0}};
   assign read_data_out_tdata[AXI4_USER_DATA_WIDTH-1:AXI4_USER_DATA_WIDTH/2] = read_data_valid_reg[1]?
      read_data_reg[FIFO_READ_DATA_UPPER_OFFSET+AXI4_CORE_DATA_WIDTH-1:FIFO_READ_DATA_UPPER_OFFSET]: {AXI4_USER_DATA_WIDTH/2{1'b0}};
   
  assign  read_data_out_tkeep[AXI4_USER_RC_TKEEP_WIDTH/2-1:0] = attr_straddle_en_i? {AXI4_USER_RC_TKEEP_WIDTH/2{1'b1}}:
      read_data_valid_reg[0]? 
      read_data_reg[AXI4_CORE_DATA_WIDTH+AXI4_CORE_RC_TKEEP_WIDTH-1:AXI4_CORE_DATA_WIDTH]: {AXI4_USER_RC_TKEEP_WIDTH/2{1'b0}};
   assign read_data_out_tkeep[AXI4_USER_RC_TKEEP_WIDTH-1:AXI4_USER_RC_TKEEP_WIDTH/2] = attr_straddle_en_i? {AXI4_USER_RC_TKEEP_WIDTH/2{1'b1}}:
      read_data_valid_reg[1]? 
      read_data_reg[FIFO_READ_TKEEP_UPPER_OFFSET+AXI4_CORE_RC_TKEEP_WIDTH-1:FIFO_READ_TKEEP_UPPER_OFFSET]:
      {AXI4_USER_RC_TKEEP_WIDTH/2{1'b0}};

   assign read_data_out_tlast = attr_straddle_en_i? 1'b0: 
      (read_data_valid_reg[0] & read_data_reg_tlast_lower) |
      (read_data_valid_reg[1] & read_data_reg_tlast_upper);

   assign output_mux_in_data = {
                read_data_out_tlast,
                read_data_out_tuser,
                read_data_out_tkeep,
                read_data_out_tdata
                };

   // Instance of output MUX
   xp4_usp_smsw_512b_rc_output_mux #
     (
      .TCQ(TCQ),
      .IMPL_TARGET(IMPL_TARGET),
      .IN_DATA_WIDTH(OUTPUT_MUX_IN_DATA_WIDTH),
      .OUT_DATA_WIDTH(AXI4_USER_DATA_WIDTH),
      .TUSER_WIDTH(AXI4_USER_RC_TUSER_WIDTH),
      .TKEEP_WIDTH(AXI4_USER_RC_TKEEP_WIDTH)
      )
     pcie_4_0_512b_rc_output_mux_blk
       (
        .clk_i(user_clk_i),
        .reset_n_i(reset_n_user_clk_i),
        .link_down_reset_i(link_down_reset_i),
    .in_data_i(output_mux_in_data),
    .in_data_valid_i(read_data_valid_reg[0]),
        .attr_straddle_en_i(attr_straddle_en_i),

    .upstream_ready_o(output_mux_ready),
    .out_data_o(m_axis_rc_tdata_o),
        .out_data_valid_o(m_axis_rc_tvalid_o),
    .out_tuser_o(m_axis_rc_tuser_o),
    .out_tlast_o(m_axis_rc_tlast_o),
    .out_tkeep_o(m_axis_rc_tkeep_o),
    .downstream_ready_i(m_axis_rc_tready_i),

    // Completion delivered indications to AXI hard block
    .pcie_compl_delivered_o(pcie_compl_delivered_user_clk),
    .pcie_compl_delivered_tag0_o(pcie_compl_delivered_tag0_user_clk),
    .pcie_compl_delivered_tag1_o(pcie_compl_delivered_tag1_user_clk),
    .pcie_compl_delivered_tag2_o(pcie_compl_delivered_tag2_user_clk),
    .pcie_compl_delivered_tag3_o(pcie_compl_delivered_tag3_user_clk)
    );

  // Return tags of delivered Completions to the AXI hard block.
  always @(posedge user_clk2_i)
    if (~reset_n_user_clk2_i)
      begin
    compl_delivered_o <= #TCQ 2'b00;
    compl_delivered_tag0_o <= #TCQ 8'd0;
    compl_delivered_tag1_o <= #TCQ 8'd0;
      end
    else if (~user_clk_en_i)
      begin
    compl_delivered_o <= #TCQ pcie_compl_delivered_user_clk[1:0];
    compl_delivered_tag0_o <= #TCQ pcie_compl_delivered_tag0_user_clk;
    compl_delivered_tag1_o <= #TCQ pcie_compl_delivered_tag1_user_clk;
      end
    else
      begin
    compl_delivered_o <= #TCQ pcie_compl_delivered_user_clk[3:2];
    compl_delivered_tag0_o <= #TCQ pcie_compl_delivered_tag2_user_clk;
    compl_delivered_tag1_o <= #TCQ pcie_compl_delivered_tag3_user_clk;
      end // else: !if(~user_clk_en_i)

endmodule // pcie_4_0_512b_rc_intfc







   
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_512b_rc_output_mux.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_512b_rc_output_mux #(
   parameter TCQ = 100,
   parameter IMPL_TARGET = "SOFT",
   parameter IN_DATA_WIDTH = 512+183+16+1,    
   parameter OUT_DATA_WIDTH = 512,
   parameter TUSER_WIDTH = 183,
   parameter TKEEP_WIDTH = 16
   )
  (
    input  wire           clk_i // 250 MHz clock for client-facing interfaces
   ,input  wire           reset_n_i // Reset in the user clock domain
   ,input  wire           link_down_reset_i // Link went down

   ,input  wire           attr_straddle_en_i // Enable straddle

   ,input wire[IN_DATA_WIDTH-1:0] in_data_i
   ,input wire in_data_valid_i
   ,output wire upstream_ready_o

   ,output reg [OUT_DATA_WIDTH-1:0]  out_data_o
   ,output reg           out_data_valid_o
   ,output reg [TUSER_WIDTH-1:0] out_tuser_o
   ,output wire          out_tlast_o
   ,output wire [TKEEP_WIDTH-1:0] out_tkeep_o
   ,input  wire           downstream_ready_i

   // Completion delivered indications to AXI hard block
   ,output reg [3:0]     pcie_compl_delivered_o
   ,output reg [7:0]     pcie_compl_delivered_tag0_o
   ,output reg [7:0]     pcie_compl_delivered_tag1_o
   ,output reg [7:0]     pcie_compl_delivered_tag2_o
   ,output reg [7:0]     pcie_compl_delivered_tag3_o
   );


   localparam MAX_CREDIT = 32;

   reg [1:0] output_fifo_occupancy;
   reg          output_fifo_write_ptr;
   reg          output_fifo_read_ptr;
   wire      output_fifo_full;
   wire      output_fifo_empty;

   reg [OUT_DATA_WIDTH-1:0] m_axis_rc_tdata_first_reg;
   reg [TKEEP_WIDTH-1:0]    m_axis_rc_tkeep_first_reg;
   reg [TUSER_WIDTH-1:0]    m_axis_rc_tuser_first_reg;
   reg                 m_axis_rc_tlast_first_reg;
   
   reg [OUT_DATA_WIDTH-1:0] m_axis_rc_tdata_second_reg;
   reg [TKEEP_WIDTH-1:0]    m_axis_rc_tkeep_second_reg;
   reg [TUSER_WIDTH-1:0]    m_axis_rc_tuser_second_reg;
   reg                 m_axis_rc_tlast_second_reg;
   
   wire             output_reg_mux_sel;
   reg                 out_tlast_reg;
   reg [TKEEP_WIDTH-1:0]    out_tkeep_reg;

  wire                 sop0_dw0;
  wire                 sop0_dw4;
  wire                 sop0_dw8;
  wire                 sop0_dw12;
  wire                 sop1_dw4;
  wire                 sop1_dw8;
  wire                 sop1_dw12;
  wire                 sop2_dw8;
  wire                 sop2_dw12;
  wire                 sop3_dw12;

   //---------------------------------------------------------------------------------------------
   // Output FIFO
   // The main FIFO feeds into two read registers in the user clock domain, which are configured
   // as a 2-entry FIFO.
   // These are termed m_axis_rc_*_reg_first and m_axis_rc_*_reg_second.
   // These can be thought of as logical extensions of the main FIFO.
   //---------------------------------------------------------------------------------------------

   // Send signal to read from main FIFO into the output FIFO when the latter is not full.
   assign    upstream_ready_o = ~output_fifo_full;

   // Maintain write and read pointers
   always @(posedge clk_i)
     if (~reset_n_i)
       output_fifo_write_ptr <= #(TCQ) 1'b0;
     else if (link_down_reset_i)
       output_fifo_write_ptr <= #(TCQ) 1'b0;
     else
       if (in_data_valid_i & ~output_fifo_full)
     output_fifo_write_ptr <= #(TCQ) ~output_fifo_write_ptr;

   always @(posedge clk_i)
     if (~reset_n_i)
       output_fifo_read_ptr <= #(TCQ) 1'b0;
     else if (link_down_reset_i)
       output_fifo_read_ptr <= #(TCQ) 1'b0;
     else
       if ((downstream_ready_i | ~out_data_valid_o) &
       ~output_fifo_empty)
     output_fifo_read_ptr <= #(TCQ) ~output_fifo_read_ptr;

    // Maintain FIFO occupancy
   always @(posedge clk_i)
     if (~reset_n_i)
       output_fifo_occupancy <= #(TCQ) 2'd0;
     else if (link_down_reset_i)
       output_fifo_occupancy <= #(TCQ) 2'd0;
     else
       if ((in_data_valid_i & ~output_fifo_full) &
       ~((downstream_ready_i | ~out_data_valid_o) &
         ~output_fifo_empty))
     output_fifo_occupancy <= #(TCQ) output_fifo_occupancy + 2'd1;
       else
     if (~(in_data_valid_i & ~output_fifo_full) &
         ((downstream_ready_i | ~out_data_valid_o) &
          ~output_fifo_empty))
       output_fifo_occupancy <= #(TCQ) output_fifo_occupancy - 2'd1;
   

   assign output_fifo_full = output_fifo_occupancy[1];
   assign output_fifo_empty = (output_fifo_occupancy == 2'b00);

   // Write data into the Output FIFO.                                                                                    
   always @(posedge clk_i)
     if (~reset_n_i)
       begin
          m_axis_rc_tdata_first_reg <= #(TCQ) {OUT_DATA_WIDTH{1'b0}};
          m_axis_rc_tdata_second_reg <= #(TCQ) {OUT_DATA_WIDTH{1'b0}};
          m_axis_rc_tkeep_first_reg <= #(TCQ) {TKEEP_WIDTH{1'b0}};
          m_axis_rc_tkeep_second_reg <= #(TCQ) {TKEEP_WIDTH{1'b0}};
          m_axis_rc_tuser_first_reg <= #(TCQ) {TUSER_WIDTH{1'b0}};
          m_axis_rc_tuser_second_reg <= #(TCQ) {TUSER_WIDTH{1'b0}};
          m_axis_rc_tlast_first_reg <= #(TCQ) 1'b0;
          m_axis_rc_tlast_second_reg <= #(TCQ) 1'b0;
       end
     else
        if (in_data_valid_i & ~output_fifo_full)
      begin
         case(output_fifo_write_ptr)
           1'b0:
         begin
            m_axis_rc_tdata_first_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH-1:0];
            m_axis_rc_tkeep_first_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH-1:OUT_DATA_WIDTH];
            m_axis_rc_tuser_first_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH+TUSER_WIDTH-1:OUT_DATA_WIDTH+TKEEP_WIDTH];
            m_axis_rc_tlast_first_reg <= #(TCQ) in_data_i[IN_DATA_WIDTH-1];
         end
           default:
         begin
            m_axis_rc_tdata_second_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH-1:0];
            m_axis_rc_tkeep_second_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH-1:OUT_DATA_WIDTH];
            m_axis_rc_tuser_second_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH+TUSER_WIDTH-1:OUT_DATA_WIDTH+TKEEP_WIDTH];
            m_axis_rc_tlast_second_reg <= #(TCQ) in_data_i[IN_DATA_WIDTH-1];
         end
         endcase // case(output_fifo_write_ptr)
      end // if (in_data_valid_i & ~output_fifo_full)
   
   // Output registers

   assign output_reg_mux_sel = output_fifo_read_ptr;

   always @(posedge clk_i)
     if (~reset_n_i)
       begin
      out_data_o <= #(TCQ) {OUT_DATA_WIDTH-1{1'b0}};
      out_tuser_o <= #(TCQ) {TUSER_WIDTH-1{1'b0}};
      out_tkeep_reg <= #(TCQ) {TKEEP_WIDTH-1{1'b0}};
      out_tlast_reg <= #(TCQ) 1'b0;
       end
     else
       if (~out_data_valid_o | downstream_ready_i)
     begin
        case(output_reg_mux_sel)
          1'b0:
        begin
           out_data_o <= #(TCQ) m_axis_rc_tdata_first_reg;
           out_tkeep_reg <= #(TCQ) m_axis_rc_tkeep_first_reg;
           out_tuser_o <= #(TCQ) m_axis_rc_tuser_first_reg;
           out_tlast_reg <= #(TCQ) m_axis_rc_tlast_first_reg;
        end
          default:
        begin
           out_data_o <= #(TCQ) m_axis_rc_tdata_second_reg;
           out_tkeep_reg <= #(TCQ) m_axis_rc_tkeep_second_reg;
           out_tuser_o <= #(TCQ) m_axis_rc_tuser_second_reg;
           out_tlast_reg <= #(TCQ) m_axis_rc_tlast_second_reg;
        end
        endcase // case(output_reg_mux_sel)
     end // if (~out_data_o | downstream_ready_i)

   always @(posedge clk_i)
     if (~reset_n_i)
       out_data_valid_o <= #(TCQ) 1'b0;
     else
       if (~out_data_valid_o | downstream_ready_i)
     out_data_valid_o <= #(TCQ) ~output_fifo_empty;

  assign out_tkeep_o =  attr_straddle_en_i? {TKEEP_WIDTH{1'b1}}: out_tkeep_reg;
  assign out_tlast_o =  attr_straddle_en_i? 1'b0: out_tlast_reg;

  //-----------------------------------------------------------------------------------------
  // Generate Completion delivered indications to AXI hard block
  //-----------------------------------------------------------------------------------------

  reg                  compl_data_valid;
  reg [3:0]          compl_delivered;
  reg              pkt_in_progress;
  reg [3:0]          compl_sop;
  reg [3:0]          compl_eop;
  reg [1:0]          compl_sop0_ptr;
  reg [1:0]          compl_sop1_ptr;
  reg [1:0]          compl_sop2_ptr;
  reg [7:0]          compl_tag0;
  reg [7:0]          compl_tag1;
  reg [7:0]          compl_tag2;
  reg [7:0]          compl_tag3;

  reg              saved_compl_delivered;
  reg [7:0]          saved_compl_tag;

  always @(posedge clk_i)
    if (~reset_n_i)
      compl_data_valid <= #(TCQ) 1'b0;
    else if (link_down_reset_i)
      compl_data_valid <= #(TCQ) 1'b0;
    else
      compl_data_valid <= #(TCQ) out_data_valid_o & downstream_ready_i;
  
  always @(posedge clk_i)
    if (~reset_n_i)
      begin
    compl_sop <= #(TCQ) 4'd0;
    compl_eop <= #(TCQ) 4'd0;
    compl_sop0_ptr <= #(TCQ) 2'd0;
    compl_sop1_ptr <= #(TCQ) 2'd0;
    compl_sop2_ptr <= #(TCQ) 2'd0;
    compl_delivered <= #(TCQ) 4'd0;
    compl_tag0 <= #(TCQ) 8'd0;
    compl_tag1 <= #(TCQ) 8'd0;
    compl_tag2 <= #(TCQ) 8'd0;
    compl_tag3 <= #(TCQ) 8'd0;
      end // if (~reset_n_i)
    else
      begin
    if (attr_straddle_en_i)
      begin
        compl_sop <= #(TCQ) out_tuser_o[67:64];
        compl_sop0_ptr <= #(TCQ) out_tuser_o[69:68];
        compl_sop1_ptr <= #(TCQ) out_tuser_o[71:70];
        compl_sop2_ptr <= #(TCQ) out_tuser_o[73:72];
        compl_eop <= #(TCQ) out_tuser_o[79:76];
        compl_delivered[0] <= #(TCQ) out_data_o[30] && (out_data_o[15:12] != 4'b0110);  // Exclude invalid tag error
        compl_delivered[1] <= #(TCQ) out_data_o[128+30] && (out_data_o[128+15:128+12] != 4'b0110);
        compl_delivered[2] <= #(TCQ) out_data_o[128*2+30] && (out_data_o[128*2+15:128*2+12] != 4'b0110);
        compl_delivered[3] <= #(TCQ) out_data_o[128*3+30] && (out_data_o[128*3+15:128*3+12] != 4'b0110);    
        compl_tag0 <= #(TCQ) out_data_o[71:64];
        compl_tag1 <= #(TCQ) out_data_o[128+71:128+64];
        compl_tag2 <= #(TCQ) out_data_o[128*2+71:128*2+64];
        compl_tag3 <= #(TCQ) out_data_o[128*3+71:128*3+64];
      end // if (attr_straddle_en_i)
    else
      begin
        compl_sop[0] <= #(TCQ) out_tuser_o[64];
        compl_sop[3:1] <= #(TCQ) 3'd0;
        compl_sop0_ptr <= #(TCQ) 2'd0;
        compl_sop1_ptr <= #(TCQ) 2'd0;
        compl_sop2_ptr <= #(TCQ) 2'd0;
        compl_eop[0] <= #(TCQ) out_tlast_reg;
        compl_eop[3:1] <= #(TCQ) 3'd0;
        compl_delivered[0] <= #(TCQ) out_data_o[30] && (out_data_o[15:12] != 4'b0110);  // Exclude invalid tag error
        compl_delivered[3:1] <= #(TCQ) 3'd0;
        compl_tag0 <= #(TCQ) out_data_o[71:64];
        compl_tag1 <= #(TCQ) 8'd0;
        compl_tag2 <= #(TCQ) 8'd0;
        compl_tag3 <= #(TCQ) 8'd0;
      end // else: !if(attr_straddle_en_i)
      end // else: !if(~reset_n_i)
    
  // Keep track of continuing packets
  always @(posedge clk_i)
    if (~reset_n_i)
      pkt_in_progress <= #(TCQ) 1'b0;
    else if (link_down_reset_i)
      pkt_in_progress <= #(TCQ) 1'b0;
    else if (compl_data_valid)
       begin
     if (attr_straddle_en_i)
       begin
         if (~pkt_in_progress)
           pkt_in_progress <= #(TCQ) ~compl_eop[0] |
                  (compl_sop[1] & ~compl_eop[1]) | 
                  (compl_sop[2] & ~compl_eop[2]) | 
                  (compl_sop[3] & ~compl_eop[3]);
         else
           pkt_in_progress <= #(TCQ) ~compl_eop[0] |
                  (compl_sop[0] & ~compl_eop[1]) | 
                  (compl_sop[1] & ~compl_eop[2]) | 
                  (compl_sop[2] & ~compl_eop[3]);
       end // if (attr_straddle_en_i)
     else
       pkt_in_progress <= #(TCQ) ~compl_eop[0];
       end // if (compl_data_valid)
    
  assign sop0_dw0 = compl_sop[0] && (compl_sop0_ptr == 2'd0) && compl_delivered[0];
  assign sop0_dw4 = compl_sop[0] && (compl_sop0_ptr == 2'd1) && compl_delivered[1];
  assign sop0_dw8 = compl_sop[0] && (compl_sop0_ptr == 2'd2) && compl_delivered[2];
  assign sop0_dw12 = compl_sop[0] && (compl_sop0_ptr == 2'd3) && compl_delivered[3];
  assign sop1_dw4 = compl_sop[1] && (compl_sop1_ptr == 2'd1) && compl_delivered[1];
  assign sop1_dw8 = compl_sop[1] && (compl_sop1_ptr == 2'd2) && compl_delivered[2];
  assign sop1_dw12 = compl_sop[1] && (compl_sop1_ptr == 2'd3) && compl_delivered[3];
  assign sop2_dw8 = compl_sop[2] && (compl_sop2_ptr == 2'd2) && compl_delivered[2];
  assign sop2_dw12 = compl_sop[2] && (compl_sop2_ptr == 2'd3) && compl_delivered[3];
  assign sop3_dw12 = compl_sop[3] & compl_delivered[3];

  // Send out tags of delivered Completions
  always @(posedge clk_i)
    if (~reset_n_i)
      begin
     pcie_compl_delivered_o <= #(TCQ) 4'd0;
     pcie_compl_delivered_tag0_o <= #(TCQ) 8'd0;
     pcie_compl_delivered_tag1_o <= #(TCQ) 8'd0;
     pcie_compl_delivered_tag2_o <= #(TCQ) 8'd0;
     pcie_compl_delivered_tag3_o <= #(TCQ) 8'd0;
      end
     else if (compl_data_valid)
       begin
     if (~pkt_in_progress)
       begin
         pcie_compl_delivered_o[0] <= #(TCQ) (sop0_dw0 & compl_eop[0])|
                      (sop1_dw4 & compl_eop[1])| 
                      (sop1_dw8 & compl_eop[1])| 
                      (sop1_dw12 & compl_eop[1])| 
                      (sop2_dw8 & compl_eop[2])| 
                      (sop2_dw12 & compl_eop[2])| 
                      (sop3_dw12 & compl_eop[3]);
         pcie_compl_delivered_tag0_o <= #(TCQ) (sop0_dw0 & compl_eop[0])?
                        compl_tag0:
                        (sop1_dw4 & compl_eop[1])? 
                        compl_tag1:
                        ((sop1_dw8 & compl_eop[1])|
                         (sop2_dw8 & compl_eop[2]))? 
                        compl_tag2:
                        compl_tag3;

         if (sop0_dw0 & compl_eop[0])
           begin
         pcie_compl_delivered_o[1] <= #(TCQ) (sop1_dw4 & compl_eop[1])| 
                          (sop1_dw8 & compl_eop[1])| 
                          (sop1_dw12 & compl_eop[1])| 
                          (sop2_dw8 & compl_eop[2])| 
                          (sop2_dw12 & compl_eop[2])| 
                          (sop3_dw12 & compl_eop[3]);
         if (sop1_dw4 & compl_eop[1])
           pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag1;
         else if ((sop1_dw8 & compl_eop[1])| 
              (sop2_dw8 & compl_eop[2]))
           pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag2;
         else
           pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag3;
           end
         else if (sop1_dw4 & compl_eop[1])
           begin
         pcie_compl_delivered_o[1] <= #(TCQ)(sop2_dw8 & compl_eop[2])| 
                          (sop2_dw12 & compl_eop[2])| 
                          (sop3_dw12 & compl_eop[3]);
         if (sop2_dw8 & compl_eop[2])
           pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag2;
         else
           pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag3;
           end
         else if (sop1_dw8 & compl_eop[1])
           begin
         pcie_compl_delivered_o[1] <= #(TCQ) sop2_dw12 & compl_eop[2];
         pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag3;
           end
         else if (sop2_dw8 & compl_eop[2])
           begin
         pcie_compl_delivered_o[1] <= #(TCQ) sop3_dw12 & compl_eop[3];
         pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag3;
           end
         else
           begin
         pcie_compl_delivered_o[1] <= #(TCQ) 1'b0;
         pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag3;
           end

         if (sop0_dw0 & compl_eop[0])
           begin
         if (sop1_dw4 & compl_eop[1])
           begin
             pcie_compl_delivered_o[2] <= #(TCQ) (sop2_dw8 & compl_eop[2])| 
                          (sop2_dw12 & compl_eop[2])| 
                          (sop3_dw12 & compl_eop[3]);
             if (sop2_dw8 & compl_eop[2])
               pcie_compl_delivered_tag2_o <= #(TCQ) compl_tag2;
             else
               pcie_compl_delivered_tag2_o <= #(TCQ) compl_tag3;
           end
         else if (sop1_dw8 & compl_eop[1])
           begin
             pcie_compl_delivered_o[2] <= #(TCQ) (sop2_dw12 & compl_eop[2])| 
                          (sop3_dw12 & compl_eop[3]);
             pcie_compl_delivered_tag2_o <= #(TCQ) compl_tag3;
           end
         else
           pcie_compl_delivered_o[2] <= #(TCQ) 1'b0;
           end // if (sop0_dw0 & compl_eop[0])
         else if (sop1_dw4 & compl_eop[1])
           begin
         if (sop2_dw8 & compl_eop[2])
           begin
             pcie_compl_delivered_o[2] <= #(TCQ) (sop3_dw12 & compl_eop[3]);
             pcie_compl_delivered_tag2_o <= #(TCQ) compl_tag3;
           end
         else
           pcie_compl_delivered_o[2] <= #(TCQ) 1'b0;
           end
         else
           pcie_compl_delivered_o[2] <= #(TCQ) 1'b0;
         
         pcie_compl_delivered_o[3] <= #(TCQ) sop0_dw0 & compl_eop[0] &
                      (sop1_dw4 & compl_eop[1]) & 
                      (sop2_dw8 & compl_eop[2]) & 
                      (sop3_dw12 & compl_eop[3]);
         pcie_compl_delivered_tag3_o <= #(TCQ) compl_tag3;
       end // if (~pkt_in_progress)
     else
       begin
         pcie_compl_delivered_o[0] <= #(TCQ) (saved_compl_delivered & compl_eop[0])|
                      (sop0_dw4 & compl_eop[1])| 
                      (sop0_dw8 & compl_eop[1])| 
                      (sop0_dw12 & compl_eop[1])| 
                      (sop1_dw8 & compl_eop[2])| 
                      (sop1_dw12 & compl_eop[2])| 
                      (sop2_dw12 & compl_eop[3]);
         pcie_compl_delivered_tag0_o <= #(TCQ) (saved_compl_delivered & compl_eop[0])?
                        saved_compl_tag:
                        (sop0_dw4 & compl_eop[1])?
                        compl_tag1:
                        ((sop0_dw8 & compl_eop[1])| 
                         (sop1_dw8 & compl_eop[2]))?
                         compl_tag2:
                         compl_tag3;

         if (saved_compl_delivered & compl_eop[0])
           begin
         pcie_compl_delivered_o[1] <= #(TCQ) (sop0_dw4 & compl_eop[1])| 
                          (sop0_dw8 & compl_eop[1])| 
                          (sop0_dw12 & compl_eop[1])| 
                          (sop1_dw8 & compl_eop[2])| 
                          (sop1_dw12 & compl_eop[2])| 
                          (sop2_dw12 & compl_eop[3]);
         if (sop0_dw4 & compl_eop[1])
           pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag1;
         else if ((sop0_dw8 & compl_eop[1])| 
              (sop1_dw8 & compl_eop[2]))
           pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag2;
         else
           pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag3;
           end
         else if (sop0_dw4 & compl_eop[1])
           begin
         pcie_compl_delivered_o[1] <= #(TCQ)(sop1_dw8 & compl_eop[2])| 
                          (sop1_dw12 & compl_eop[2])| 
                          (sop2_dw12 & compl_eop[3]);
         if (sop1_dw8 & compl_eop[2])
           pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag2;
         else
           pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag3;
           end
         else if (sop0_dw8 & compl_eop[1])
           begin
         pcie_compl_delivered_o[1] <= #(TCQ) sop1_dw12 & compl_eop[2];
         pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag3;
           end
         else if (sop1_dw8 & compl_eop[2])
           begin
         pcie_compl_delivered_o[1] <= #(TCQ) sop2_dw12 & compl_eop[3];
         pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag3;
           end
         else
           begin
         pcie_compl_delivered_o[1] <= #(TCQ) 1'b0;
         pcie_compl_delivered_tag1_o <= #(TCQ) compl_tag3;
           end

         if (saved_compl_delivered & compl_eop[0])
           begin
         if (sop0_dw4 & compl_eop[1])
           begin
             pcie_compl_delivered_o[2] <= #(TCQ) (sop1_dw8 & compl_eop[2])| 
                          (sop1_dw12 & compl_eop[2])| 
                          (sop2_dw12 & compl_eop[3]);
             if (sop1_dw8 & compl_eop[2])
               pcie_compl_delivered_tag2_o <= #(TCQ) compl_tag2;
             else
               pcie_compl_delivered_tag2_o <= #(TCQ) compl_tag3;
           end
         else if (sop0_dw8 & compl_eop[1])
           begin
             pcie_compl_delivered_o[2] <= #(TCQ) (sop1_dw12 & compl_eop[2])| 
                          (sop2_dw12 & compl_eop[3]);
             pcie_compl_delivered_tag2_o <= #(TCQ) compl_tag3;
           end
         else
           pcie_compl_delivered_o[2] <= #(TCQ) 1'b0;
           end // if (saved_compl_delivered & compl_eop[0])
         else if (sop0_dw4 & compl_eop[1])
           begin
         if (sop1_dw8 & compl_eop[2])
           begin
             pcie_compl_delivered_o[2] <= #(TCQ) (sop2_dw12 & compl_eop[3]);
             pcie_compl_delivered_tag2_o <= #(TCQ) compl_tag3;
           end
         else
           pcie_compl_delivered_o[2] <= #(TCQ) 1'b0;
           end
         else
           pcie_compl_delivered_o[2] <= #(TCQ) 1'b0;

         pcie_compl_delivered_o[3] <= #(TCQ) (saved_compl_delivered & compl_eop[0]) &
                      (sop0_dw4 & compl_eop[1]) & 
                      (sop1_dw8 & compl_eop[2]) & 
                      (sop2_dw12 & compl_eop[3]);
         pcie_compl_delivered_tag3_o <= #(TCQ) compl_tag3;
       end // else: !if(~pkt_in_progress)
       end // if (compl_data_valid)
     else
       pcie_compl_delivered_o <= #(TCQ) 4'd0;

  // Save tag for next cycle
   always @(posedge clk_i)
     if (~reset_n_i)
       begin
     saved_compl_delivered <= #(TCQ) 1'b0;
     saved_compl_tag <= #(TCQ) 8'd0;
       end
     else if (compl_data_valid)
       begin
     if (compl_sop[3])
       begin
         saved_compl_delivered <= #(TCQ) compl_delivered[3];
         saved_compl_tag <= #(TCQ) compl_tag3;
       end
     else if (compl_sop[2])
       case(compl_sop2_ptr)
         2'd2:
           begin
         saved_compl_delivered <= #(TCQ) compl_delivered[2];
         saved_compl_tag <= #(TCQ) compl_tag2;
           end
         default:
           begin
         saved_compl_delivered <= #(TCQ) compl_delivered[3];
         saved_compl_tag <= #(TCQ) compl_tag3;
           end
       endcase // case(compl_sop2_ptr)
     else if (compl_sop[1])
       case(compl_sop1_ptr)
         2'd1:
           begin
         saved_compl_delivered <= #(TCQ) compl_delivered[1];
         saved_compl_tag <= #(TCQ) compl_tag1;
           end
         2'd2:
           begin
         saved_compl_delivered <= #(TCQ) compl_delivered[2];
         saved_compl_tag <= #(TCQ) compl_tag2;
           end
         default:
           begin
         saved_compl_delivered <= #(TCQ) compl_delivered[3];
         saved_compl_tag <= #(TCQ) compl_tag3;
           end
       endcase // case(compl_sop1_ptr)
     else if (compl_sop[0])
       case(compl_sop0_ptr)
         2'd0:
           begin
         saved_compl_delivered <= #(TCQ) compl_delivered[0];
         saved_compl_tag <= #(TCQ) compl_tag0;
           end
         2'd1:
           begin
         saved_compl_delivered <= #(TCQ) compl_delivered[1];
         saved_compl_tag <= #(TCQ) compl_tag1;
           end
         2'd2:
           begin
         saved_compl_delivered <= #(TCQ) compl_delivered[2];
         saved_compl_tag <= #(TCQ) compl_tag2;
           end
         default:
           begin
         saved_compl_delivered <= #(TCQ) compl_delivered[3];
         saved_compl_tag <= #(TCQ) compl_tag3;
           end
       endcase // case(compl_sop0_ptr)
       end // if (compl_data_valid)

endmodule // pcie_4_0_512b_rc_output_mux
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_512b_rq_intfc.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_512b_rq_intfc #(
   parameter TCQ = 100,
   parameter IMPL_TARGET = "SOFT",
   parameter AXI4_USER_DATA_WIDTH = 512,
   parameter AXI4_CORE_DATA_WIDTH = 256,
   parameter AXI4_USER_RQ_TUSER_WIDTH = 137,
   parameter AXI4_CORE_RQ_TUSER_WIDTH = 62,
   parameter AXI4_USER_RQ_TKEEP_WIDTH = 16,
   parameter AXI4_CORE_RQ_TKEEP_WIDTH = 8,
   parameter AXI4_CORE_RQ_TREADY_WIDTH = 4,
   parameter PARITY_ENABLE = 0                
   ) 
  (
    input  wire           user_clk2_i // 500 MHz clock for core-facing interfaces
   ,input  wire           user_clk_i // 250 MHz clock for client-facing interfaces
   ,input  wire           user_clk_en_i // User clock enable for clock domain crossing
   ,input  wire           reset_n_user_clk_i // Reset in the user clock domain
   ,input  wire           reset_n_user_clk2_i // Reset in the user clock2 domain
   ,input  wire           link_down_reset_i // Link went down
   // Attributes
   ,input  wire           attr_straddle_en_i // Enable straddle
   ,input wire [1:0]      attr_alignment_mode_i // Payload alignment mode
                                                // (00= Dword-aligned, 10 = 128b address-aligned)
   ,input wire            attr_axisten_if_rq_cc_registered_tready_i // 0 = registered_tready enabled, 1 = registered_tready disabled
   //-----------------------------------------------------------------------------------------------
   // Client-side signals
   //-----------------------------------------------------------------------------------------------
   ,input wire [511:0]    s_axis_rq_tdata_i
   ,input wire            s_axis_rq_tvalid_i
   ,input wire [AXI4_USER_RQ_TUSER_WIDTH-1:0] s_axis_rq_tuser_i
   ,input wire            s_axis_rq_tlast_i
   ,input wire [AXI4_USER_RQ_TKEEP_WIDTH-1:0] s_axis_rq_tkeep_i
   ,output reg            s_axis_rq_tready_o   
   //-----------------------------------------------------------------------------------------------
   // Core-side signals
   //-----------------------------------------------------------------------------------------------
   ,output wire [255:0]   core_rq_tdata_o
   ,output wire           core_rq_tvalid_o
   ,output wire [AXI4_CORE_RQ_TUSER_WIDTH-1:0] core_rq_tuser_o
   ,output wire            core_rq_tlast_o
   ,output wire [AXI4_CORE_RQ_TKEEP_WIDTH-1:0] core_rq_tkeep_o
   ,input wire [AXI4_CORE_RQ_TREADY_WIDTH-1:0] core_rq_tready_i
   );

   localparam FIFO_IN_DATA_WIDTH = AXI4_USER_DATA_WIDTH + AXI4_USER_RQ_TKEEP_WIDTH + AXI4_CORE_RQ_TUSER_WIDTH*2 +
                   2; // tlast
   localparam FIFO_OUT_DATA_WIDTH = FIFO_IN_DATA_WIDTH/2;

   localparam OUTPUT_MUX_IN_DATA_WIDTH = AXI4_CORE_DATA_WIDTH + AXI4_CORE_RQ_TKEEP_WIDTH + AXI4_CORE_RQ_TUSER_WIDTH + 1;

   reg [AXI4_USER_DATA_WIDTH-1:0] s_axis_rq_tdata_reg;
   reg                   s_axis_rq_tvalid_reg_lower;
   reg                   s_axis_rq_tvalid_reg_upper;
   reg [AXI4_USER_RQ_TKEEP_WIDTH-1:0] s_axis_rq_tkeep_reg;
   reg                       s_axis_rq_tlast_reg_lower;
   reg                       s_axis_rq_tlast_reg_upper;
   reg [AXI4_USER_RQ_TUSER_WIDTH-1:0] s_axis_rq_tuser_reg;


   wire [1:0]                   s_axis_rq_sop;
   wire [1:0]                   s_axis_rq_eop;
   wire [1:0]                   s_axis_rq_sop0_ptr;
   wire [3:0]                   s_axis_rq_eop0_ptr;
   wire [3:0]                   s_axis_rq_eop1_ptr;
   wire [63:0]                   s_axis_rq_parity;

   wire [AXI4_CORE_RQ_TUSER_WIDTH*2-1:0] fifo_in_data_tuser;
   wire [1:0]                  fifo_in_data_tlast;

   wire [FIFO_IN_DATA_WIDTH-1:0]      fifo_in_data;
   wire [1:0]                  fifo_in_data_valid;
   wire                  fifo_almost_full_user_clk;

   reg                      s_axis_rq_tuser_discontinue_reg_lower;
   reg                      s_axis_rq_tuser_discontinue_reg_upper;

    wire [FIFO_OUT_DATA_WIDTH-1:0]      fifo_read_data;
   wire                  fifo_read_data_valid;
   wire                  output_mux_ready;

  wire [3:0] 		 s_axis_rq_fbe_lower;
  wire [3:0] 		 s_axis_rq_fbe_upper;
  wire [3:0] 		 s_axis_rq_lbe_lower;
  wire [3:0] 		 s_axis_rq_lbe_upper;
  wire [1:0]             s_axis_rq_addr_offset_lower;
  wire [1:0]             s_axis_rq_addr_offset_upper;
  wire 			 s_axis_rq_tph_present_lower;
  wire 			 s_axis_rq_tph_present_upper;
  wire [1:0] 		 s_axis_rq_tph_type_lower;
  wire [1:0] 		 s_axis_rq_tph_type_upper;
  wire [7:0] 		 s_axis_rq_tph_st_tag_lower;
  wire [7:0] 		 s_axis_rq_tph_st_tag_upper;
  wire [5:0] 		 s_axis_rq_seq_num_lower;
  wire [5:0] 		 s_axis_rq_seq_num_upper;
  wire [63:0] 		 s_axis_rq_parity_i;

  reg [AXI4_CORE_RQ_TREADY_WIDTH-1:0] core_rq_tready_reg;
  wire [AXI4_CORE_RQ_TREADY_WIDTH-1:0] core_rq_tready_int;

  assign  s_axis_rq_sop[1:0] =  s_axis_rq_tuser_i[21:20];
  assign  s_axis_rq_sop0_ptr[1:0] =  s_axis_rq_tuser_i[23:22];
  assign  s_axis_rq_eop[1:0] =  s_axis_rq_tuser_i[27:26];
  assign  s_axis_rq_eop0_ptr[3:0] =  s_axis_rq_tuser_i[31:28];
  assign  s_axis_rq_eop1_ptr[3:0] =  s_axis_rq_tuser_i[35:32];

  // First BE
  assign  s_axis_rq_fbe_lower[3:0] = s_axis_rq_tuser_i[3:0];
  assign  s_axis_rq_fbe_upper[3:0] = (attr_straddle_en_i & s_axis_rq_sop[0] & s_axis_rq_sop0_ptr[1])?
	  s_axis_rq_tuser_i[3:0]: s_axis_rq_tuser_i[7:4];
  // Last BE
  assign  s_axis_rq_lbe_lower[3:0] = s_axis_rq_tuser_i[11:8];
  assign  s_axis_rq_lbe_upper[3:0] =  (attr_straddle_en_i & s_axis_rq_sop[0] & s_axis_rq_sop0_ptr[1])? 
	  s_axis_rq_tuser_i[11:8]: s_axis_rq_tuser_i[15:12];
  // Address Offset
  assign  s_axis_rq_addr_offset_lower[1:0] = s_axis_rq_tuser_i[17:16];
  assign  s_axis_rq_addr_offset_upper[1:0] = (attr_straddle_en_i & s_axis_rq_sop[0] & s_axis_rq_sop0_ptr[1])?
	  s_axis_rq_tuser_i[17:16]: s_axis_rq_tuser_i[19:18];
  // TPH-related signals
  assign  s_axis_rq_tph_present_lower = s_axis_rq_tuser_i[37];
  assign  s_axis_rq_tph_present_upper = (attr_straddle_en_i & s_axis_rq_sop[0] & s_axis_rq_sop0_ptr[1])?
	  s_axis_rq_tuser_i[37]: s_axis_rq_tuser_i[38];
  assign  s_axis_rq_tph_type_lower[1:0] = s_axis_rq_tuser_i[40:39];
  assign  s_axis_rq_tph_type_upper[1:0] = (attr_straddle_en_i & s_axis_rq_sop[0] & s_axis_rq_sop0_ptr[1])?
	  s_axis_rq_tuser_i[40:39]: s_axis_rq_tuser_i[42:41];
  assign  s_axis_rq_tph_st_tag_lower[7:0] = s_axis_rq_tuser_i[52:45];
  assign  s_axis_rq_tph_st_tag_upper[7:0] = (attr_straddle_en_i & s_axis_rq_sop[0] & s_axis_rq_sop0_ptr[1])?
	  s_axis_rq_tuser_i[52:45]: s_axis_rq_tuser_i[60:53];
  assign  s_axis_rq_seq_num_lower[5:0] = s_axis_rq_tuser_i[66:61];
  assign  s_axis_rq_seq_num_upper[5:0] = (attr_straddle_en_i & s_axis_rq_sop[0] & s_axis_rq_sop0_ptr[1])?
	  s_axis_rq_tuser_i[66:61]: s_axis_rq_tuser_i[72:67];
  // Parity
  generate
    if (PARITY_ENABLE)
      assign  s_axis_rq_parity_i[63:0] =  s_axis_rq_tuser_i[136:73];
    else
      assign  s_axis_rq_parity_i[63:0] =  64'd0;
  endgenerate    

   // Register input data
   always @(posedge user_clk_i)
     if (~reset_n_user_clk_i)
       begin
      s_axis_rq_tdata_reg <= {AXI4_USER_DATA_WIDTH{1'b0}};
      s_axis_rq_tvalid_reg_lower <= 1'b0;
      s_axis_rq_tvalid_reg_upper <= 1'b0;
      s_axis_rq_tkeep_reg <= {AXI4_USER_RQ_TKEEP_WIDTH{1'b0}};
      s_axis_rq_tuser_reg <= {AXI4_USER_RQ_TUSER_WIDTH{1'b0}};
      s_axis_rq_tuser_discontinue_reg_lower <= 1'b0;
       s_axis_rq_tuser_discontinue_reg_upper <= 1'b0;
      s_axis_rq_tlast_reg_lower <= 1'b0;
      s_axis_rq_tlast_reg_upper <= 1'b0;
       end
     else
       begin
      s_axis_rq_tdata_reg <= s_axis_rq_tdata_i;
      s_axis_rq_tvalid_reg_lower <= s_axis_rq_tvalid_i & s_axis_rq_tready_o;
      s_axis_rq_tvalid_reg_upper <= attr_straddle_en_i? (~s_axis_rq_eop[0] | s_axis_rq_eop0_ptr[3] |
                                 (s_axis_rq_sop[0] & s_axis_rq_sop0_ptr[1]) |
                                 s_axis_rq_sop[1]) &
                    s_axis_rq_tvalid_i & s_axis_rq_tready_o:
                    (~s_axis_rq_tlast_i | s_axis_rq_tkeep_i[8]) &
                    s_axis_rq_tvalid_i & s_axis_rq_tready_o;
     // Generate tkeep settings for core side
     if (~attr_straddle_en_i)
       s_axis_rq_tkeep_reg[7:0] <= s_axis_rq_tkeep_i[7:0];
     else if (s_axis_rq_tvalid_i & s_axis_rq_tready_o)
       begin
         if (~s_axis_rq_eop[0] | s_axis_rq_eop0_ptr[3])
           s_axis_rq_tkeep_reg[7:0] <= 8'hff;
         else
           case(s_axis_rq_eop0_ptr[2:0])
         3'd0: s_axis_rq_tkeep_reg[7:0] <= 8'h01;
         3'd1: s_axis_rq_tkeep_reg[7:0] <= 8'h03;
         3'd2: s_axis_rq_tkeep_reg[7:0] <= 8'h07;
         3'd3: s_axis_rq_tkeep_reg[7:0] <= 8'h0f;
         3'd4: s_axis_rq_tkeep_reg[7:0] <= 8'h1f;
         3'd5: s_axis_rq_tkeep_reg[7:0] <= 8'h3f;
         3'd6: s_axis_rq_tkeep_reg[7:0] <= 8'h7f;
         default: s_axis_rq_tkeep_reg[7:0] <= 8'hff;
           endcase // case(s_axis_rq_eop0_ptr[2:0])
       end // if (s_axis_rq_tvalid_i & s_axis_rq_tready_o)
     else
       s_axis_rq_tkeep_reg[7:0] <= 8'd0;
         
     if (~attr_straddle_en_i)
       s_axis_rq_tkeep_reg[15:8] <= s_axis_rq_tkeep_i[15:8];
     else if (s_axis_rq_tvalid_i & s_axis_rq_tready_o)
       begin
         if (~s_axis_rq_eop[0])
           s_axis_rq_tkeep_reg[15:8] <= 8'hff;
         else if (s_axis_rq_eop0_ptr[3])
           case(s_axis_rq_eop0_ptr[2:0])
         3'd0: s_axis_rq_tkeep_reg[15:8] <= 8'h01;
         3'd1: s_axis_rq_tkeep_reg[15:8] <= 8'h03;
         3'd2: s_axis_rq_tkeep_reg[15:8] <= 8'h07;
         3'd3: s_axis_rq_tkeep_reg[15:8] <= 8'h0f;
         3'd4: s_axis_rq_tkeep_reg[15:8] <= 8'h1f;
         3'd5: s_axis_rq_tkeep_reg[15:8] <= 8'h3f;
         3'd6: s_axis_rq_tkeep_reg[15:8] <= 8'h7f;
         default: s_axis_rq_tkeep_reg[15:8] <= 8'hff;
           endcase // case(s_axis_rq_eop0_ptr[2:0])
         else if ((s_axis_rq_sop[0] && (s_axis_rq_sop0_ptr[1]))||
              s_axis_rq_sop[1])
           // Packet starting in second half
           begin
         if (~s_axis_rq_eop[1])
           s_axis_rq_tkeep_reg[15:8] <= 8'hff;
         else
           case(s_axis_rq_eop1_ptr[2:0])
             3'd2: s_axis_rq_tkeep_reg[15:8] <= 8'h07;
             3'd3: s_axis_rq_tkeep_reg[15:8] <= 8'h0f;
             3'd4: s_axis_rq_tkeep_reg[15:8] <= 8'h1f;
             3'd5: s_axis_rq_tkeep_reg[15:8] <= 8'h3f;
             3'd6: s_axis_rq_tkeep_reg[15:8] <= 8'h7f;
             default: s_axis_rq_tkeep_reg[15:8] <= 8'hff;
           endcase // case(s_axis_rq_eop1_ptr[2:0])
           end // if ((s_axis_rq_sop[0] && (s_axis_rq_sop0_ptr[1]))||...
         else
           s_axis_rq_tkeep_reg[15:8] <= 8'd0;
       end // if (s_axis_rq_tvalid_i & s_axis_rq_tready_o)
     else
       s_axis_rq_tkeep_reg[15:8] <= 8'd0;


      s_axis_rq_tuser_reg <= {
			      s_axis_rq_parity_i[63:0],
			      s_axis_rq_seq_num_upper[5:0],
			      s_axis_rq_seq_num_lower[5:0],
			      s_axis_rq_tph_st_tag_upper[7:0],
			      s_axis_rq_tph_st_tag_lower[7:0],
			      2'd0, // TPH Indirect Tag Enable
			      s_axis_rq_tph_type_upper[1:0],
			      s_axis_rq_tph_type_lower[1:0],
			      s_axis_rq_tph_present_upper,
			      s_axis_rq_tph_present_lower,
			      s_axis_rq_tuser_i[36:20],
			      s_axis_rq_addr_offset_upper[1:0],
			      s_axis_rq_addr_offset_lower[1:0],
			      s_axis_rq_lbe_upper[3:0],
			      s_axis_rq_lbe_lower[3:0],
			      s_axis_rq_fbe_upper[3:0],
			      s_axis_rq_fbe_lower[3:0]
			      };

     // Generate discontinue for lower and upper halves
     if (~attr_straddle_en_i) 
       begin
         s_axis_rq_tuser_discontinue_reg_lower <= s_axis_rq_tuser_i[36] &
                              (~s_axis_rq_tlast_i |
                               ~s_axis_rq_tkeep_i[8]);
         s_axis_rq_tuser_discontinue_reg_upper <= s_axis_rq_tuser_i[36] &
                              (~s_axis_rq_tlast_i |
                               s_axis_rq_tkeep_i[8]);
       end // if (~attr_straddle_en_i)
     else
       begin
         s_axis_rq_tuser_discontinue_reg_lower <= s_axis_rq_tuser_i[36] &
                              (~s_axis_rq_eop[0] |
                               ~s_axis_rq_eop0_ptr[3]);
         s_axis_rq_tuser_discontinue_reg_upper <= s_axis_rq_tuser_i[36] &
                              (~s_axis_rq_eop[0] |
                               s_axis_rq_eop0_ptr[3]);
       end // else: !if(~attr_straddle_en_i)
     
     s_axis_rq_tlast_reg_lower <= attr_straddle_en_i? 
                      (s_axis_rq_eop[0] & ~s_axis_rq_eop0_ptr[3]):
                      (s_axis_rq_tlast_i & ~s_axis_rq_tkeep_i[8]);
     s_axis_rq_tlast_reg_upper <= attr_straddle_en_i? 
                      (s_axis_rq_eop[0] & s_axis_rq_eop0_ptr[3]) | s_axis_rq_eop[1]:
                      (s_axis_rq_tlast_i & s_axis_rq_tkeep_i[8]);
       end // else: !if(~reset_n_user_clk_i)

  assign s_axis_rq_parity[63:0] =  PARITY_ENABLE? s_axis_rq_tuser_reg[136:73] : 64'd0;

   // Generate the tuser signals for the core side
   // discontinue
  assign  fifo_in_data_tuser[11] = s_axis_rq_tuser_discontinue_reg_lower;
   assign fifo_in_data_tuser[AXI4_CORE_RQ_TUSER_WIDTH+11] = s_axis_rq_tuser_discontinue_reg_upper;

  // First and Last BE
  assign  fifo_in_data_tuser[3:0] = s_axis_rq_tuser_reg[3:0]; // First BE
  assign  fifo_in_data_tuser[AXI4_CORE_RQ_TUSER_WIDTH+3:AXI4_CORE_RQ_TUSER_WIDTH] = s_axis_rq_tuser_reg[7:4];
  assign  fifo_in_data_tuser[7:4] = s_axis_rq_tuser_reg[11:8]; // Last BE
  assign  fifo_in_data_tuser[AXI4_CORE_RQ_TUSER_WIDTH+7:AXI4_CORE_RQ_TUSER_WIDTH+4] = s_axis_rq_tuser_reg[15:12];

  // addr offset
  assign  fifo_in_data_tuser[10:8] = {1'b0, s_axis_rq_tuser_reg[17:16]}; 
  assign  fifo_in_data_tuser[AXI4_CORE_RQ_TUSER_WIDTH+10:AXI4_CORE_RQ_TUSER_WIDTH+8] =
      {1'b0, s_axis_rq_tuser_reg[19:18]}; 
  // TPH present
  assign  fifo_in_data_tuser[12] = s_axis_rq_tuser_reg[37];
  assign  fifo_in_data_tuser[AXI4_CORE_RQ_TUSER_WIDTH+12] =s_axis_rq_tuser_reg[38];
  // TPH Type
  assign  fifo_in_data_tuser[14:13] = s_axis_rq_tuser_reg[40:39];
  assign  fifo_in_data_tuser[AXI4_CORE_RQ_TUSER_WIDTH+14:AXI4_CORE_RQ_TUSER_WIDTH+13] = s_axis_rq_tuser_reg[42:41];
  // TPH Indirect Tag Enable
  assign  fifo_in_data_tuser[15] = 1'b0;
  assign  fifo_in_data_tuser[AXI4_CORE_RQ_TUSER_WIDTH+15] = 1'b0;
  // TPH Steering Tag
  assign  fifo_in_data_tuser[23:16] = s_axis_rq_tuser_reg[52:45];
  assign  fifo_in_data_tuser[AXI4_CORE_RQ_TUSER_WIDTH+23:AXI4_CORE_RQ_TUSER_WIDTH+16] = s_axis_rq_tuser_reg[60:53];
  // Sequence Number
  assign  fifo_in_data_tuser[27:24] = s_axis_rq_tuser_reg[64:61];
  assign  fifo_in_data_tuser[61:60] = s_axis_rq_tuser_reg[66:65];
  assign  fifo_in_data_tuser[AXI4_CORE_RQ_TUSER_WIDTH+27:AXI4_CORE_RQ_TUSER_WIDTH+24] = s_axis_rq_tuser_reg[70:67];
  assign  fifo_in_data_tuser[AXI4_CORE_RQ_TUSER_WIDTH+61:AXI4_CORE_RQ_TUSER_WIDTH+60] = s_axis_rq_tuser_reg[72:71];
   // parity
   assign fifo_in_data_tuser[59:28] = s_axis_rq_parity[31:0];
   assign fifo_in_data_tuser[AXI4_CORE_RQ_TUSER_WIDTH+59:AXI4_CORE_RQ_TUSER_WIDTH+28] = s_axis_rq_parity[63:32];
   
   // Generate tlast for lower and upper halves
  assign fifo_in_data_tlast[0] = s_axis_rq_tlast_reg_lower;
  assign fifo_in_data_tlast[1] = s_axis_rq_tlast_reg_upper;

   // Generate valid for upper half
  assign fifo_in_data_valid[0] = s_axis_rq_tvalid_reg_lower;
  assign fifo_in_data_valid[1] = s_axis_rq_tvalid_reg_upper;

   assign fifo_in_data[AXI4_CORE_DATA_WIDTH-1:0] = s_axis_rq_tdata_reg[AXI4_CORE_DATA_WIDTH-1:0];
   assign fifo_in_data[FIFO_IN_DATA_WIDTH/2+AXI4_CORE_DATA_WIDTH-1:FIFO_IN_DATA_WIDTH/2] =
      s_axis_rq_tdata_reg[AXI4_CORE_DATA_WIDTH*2-1:AXI4_CORE_DATA_WIDTH];

   assign fifo_in_data[AXI4_CORE_DATA_WIDTH + AXI4_CORE_RQ_TKEEP_WIDTH-1: AXI4_CORE_DATA_WIDTH] =
      s_axis_rq_tkeep_reg[AXI4_CORE_RQ_TKEEP_WIDTH-1:0];
  assign  fifo_in_data[FIFO_IN_DATA_WIDTH/2 + AXI4_CORE_DATA_WIDTH + AXI4_CORE_RQ_TKEEP_WIDTH-1:
               FIFO_IN_DATA_WIDTH/2 + AXI4_CORE_DATA_WIDTH] =
      s_axis_rq_tkeep_reg[AXI4_CORE_RQ_TKEEP_WIDTH*2-1:AXI4_CORE_RQ_TKEEP_WIDTH];

   assign fifo_in_data[AXI4_CORE_DATA_WIDTH + AXI4_CORE_RQ_TKEEP_WIDTH +  AXI4_CORE_RQ_TUSER_WIDTH-1:
               AXI4_CORE_DATA_WIDTH + AXI4_CORE_RQ_TKEEP_WIDTH] = 
      fifo_in_data_tuser[AXI4_CORE_RQ_TUSER_WIDTH-1:0];
   assign fifo_in_data[FIFO_IN_DATA_WIDTH/2 + AXI4_CORE_DATA_WIDTH + AXI4_CORE_RQ_TKEEP_WIDTH +  AXI4_CORE_RQ_TUSER_WIDTH-1:
               FIFO_IN_DATA_WIDTH/2 + AXI4_CORE_DATA_WIDTH + AXI4_CORE_RQ_TKEEP_WIDTH] = 
      fifo_in_data_tuser[AXI4_CORE_RQ_TUSER_WIDTH*2-1:AXI4_CORE_RQ_TUSER_WIDTH];

   assign fifo_in_data[AXI4_CORE_DATA_WIDTH + AXI4_CORE_RQ_TKEEP_WIDTH +  AXI4_CORE_RQ_TUSER_WIDTH] =
      fifo_in_data_tlast[0];
   assign fifo_in_data[FIFO_IN_DATA_WIDTH/2 + AXI4_CORE_DATA_WIDTH + AXI4_CORE_RQ_TKEEP_WIDTH +  AXI4_CORE_RQ_TUSER_WIDTH] =
      fifo_in_data_tlast[1];
 
   // De-assert ready when FIFO is almost full
   always @(posedge user_clk_i)
     if (~reset_n_user_clk_i)
       s_axis_rq_tready_o <= 1'b0;
     else
       s_axis_rq_tready_o <= #(TCQ) ~fifo_almost_full_user_clk;

  // Register tready from hard block
   always @(posedge user_clk2_i)
     if (~reset_n_user_clk2_i)
       core_rq_tready_reg <= {AXI4_CORE_RQ_TREADY_WIDTH{1'b0}};
     else
       core_rq_tready_reg <= core_rq_tready_i;

  assign  core_rq_tready_int = attr_axisten_if_rq_cc_registered_tready_i?
      core_rq_tready_reg : core_rq_tready_i;

   // Async FIFO
   xp4_usp_smsw_512b_async_fifo #
     (
      .TCQ(TCQ),
      .IMPL_TARGET(IMPL_TARGET),
      .IN_DATA_WIDTH(FIFO_IN_DATA_WIDTH),
      .FIFO_WIDTH(FIFO_OUT_DATA_WIDTH),
      .FIFO_DEPTH(16),
      .FIFO_ALMOST_FULL_THRESHOLD(7)
      )
     pcie_4_0_512b_async_fifo_blk
       (
    .clk_i(user_clk2_i),
    .clk_en_i(user_clk_en_i),
        .reset_n_i(reset_n_user_clk2_i),
        .link_down_reset_i(link_down_reset_i),
    // Write side
    .write_data_i(fifo_in_data),
    .write_en_i(fifo_in_data_valid),
    .fifo_almost_full_o(fifo_almost_full_user_clk),
    // Read side
    .read_en_i(output_mux_ready),
    .read_data_o(fifo_read_data),
    .read_data_valid_o(fifo_read_data_valid)
    );

   // Instance of output MUX
   xp4_usp_smsw_512b_rq_output_mux #
     (
      .TCQ(TCQ),
      .IMPL_TARGET(IMPL_TARGET),
      .IN_DATA_WIDTH(OUTPUT_MUX_IN_DATA_WIDTH),
      .OUT_DATA_WIDTH(AXI4_CORE_DATA_WIDTH),
      .TUSER_WIDTH(AXI4_CORE_RQ_TUSER_WIDTH),
      .TKEEP_WIDTH(AXI4_CORE_RQ_TKEEP_WIDTH),
      .TREADY_WIDTH(AXI4_CORE_RQ_TREADY_WIDTH)
      )
     pcie_4_0_512b_rq_output_mux_blk
       (
        .clk_i(user_clk2_i),
        .reset_n_i(reset_n_user_clk_i),
        .link_down_reset_i(link_down_reset_i),
    .in_data_i(fifo_read_data),
    .in_data_valid_i(fifo_read_data_valid),
    .upstream_ready_o(output_mux_ready),

    .out_data_o(core_rq_tdata_o),
        .out_data_valid_o(core_rq_tvalid_o),
    .out_tuser_o(core_rq_tuser_o),
    .out_tlast_o(core_rq_tlast_o),
    .out_tkeep_o(core_rq_tkeep_o),
    .downstream_ready_i(core_rq_tready_int)
    );

endmodule // pcie_4_0_512b_rq_intfc







   
//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_512b_rq_output_mux.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_512b_rq_output_mux #(
   parameter TCQ = 100,
   parameter IMPL_TARGET = "SOFT",
   parameter IN_DATA_WIDTH = 256+33+8+1,    
   parameter OUT_DATA_WIDTH = 256,
   parameter TUSER_WIDTH = 33,
   parameter TKEEP_WIDTH = 8,
   parameter TREADY_WIDTH = 4
   )
  (
    input  wire           clk_i // 250 MHz clock for client-facing interfaces
   ,input  wire           reset_n_i // Reset in the user clock domain
   ,input  wire           link_down_reset_i // Link went down

   ,input wire[IN_DATA_WIDTH-1:0] in_data_i
   ,input wire in_data_valid_i
   ,output wire upstream_ready_o

   ,output reg [OUT_DATA_WIDTH-1:0]  out_data_o
   ,output reg           out_data_valid_o
   ,output reg [TUSER_WIDTH-1:0] out_tuser_o
   ,output reg          out_tlast_o
   ,output reg [TKEEP_WIDTH-1:0] out_tkeep_o
   ,input  wire [TREADY_WIDTH-1:0]  downstream_ready_i
   );


   reg [1:0] output_fifo_occupancy;
  reg          output_fifo_write_ptr;
  reg          output_fifo_read_ptr;
   wire      output_fifo_full;
   wire      output_fifo_empty;

   reg [OUT_DATA_WIDTH-1:0] m_axis_rq_tdata_first_reg;
   reg [TKEEP_WIDTH-1:0]    m_axis_rq_tkeep_first_reg;
   reg [TUSER_WIDTH-1:0]    m_axis_rq_tuser_first_reg;
   reg                 m_axis_rq_tlast_first_reg;
   
   reg [OUT_DATA_WIDTH-1:0] m_axis_rq_tdata_second_reg;
   reg [TKEEP_WIDTH-1:0]    m_axis_rq_tkeep_second_reg;
   reg [TUSER_WIDTH-1:0]    m_axis_rq_tuser_second_reg;
   reg                 m_axis_rq_tlast_second_reg;
   
   wire             output_reg_mux_sel;
   //---------------------------------------------------------------------------------------------
   // Output FIFO.
   // The main FIFO feeds into two read registers in the core clock domain, which are configured
   // as a 2-entry FIFO.
   // This can be thought of as logical extensions of the main FIFO.
   //---------------------------------------------------------------------------------------------

   assign    upstream_ready_o = ~output_fifo_full;

   // Maintain write and read pointers
   // Write pointer is updated only in alternate cycles.
   always @(posedge clk_i)
     if (~reset_n_i)
       output_fifo_write_ptr <= #(TCQ)  1'b0;
     else if (link_down_reset_i)
       output_fifo_write_ptr <= #(TCQ)  1'b0;
     else
       if (in_data_valid_i & ~output_fifo_full)
     output_fifo_write_ptr <= #(TCQ) ~output_fifo_write_ptr;
   
   always @(posedge clk_i)
     if (~reset_n_i)
       output_fifo_read_ptr <= #(TCQ) 2'd0;
     else if (link_down_reset_i)
       output_fifo_read_ptr <= #(TCQ) 2'd0;
     else
       if ((downstream_ready_i[3] | ~out_data_valid_o) &
       ~output_fifo_empty)
     output_fifo_read_ptr <= #(TCQ) ~output_fifo_read_ptr;

      // Maintain FIFO occupancy
   always @(posedge clk_i)
     if (~reset_n_i)
       output_fifo_occupancy <= #(TCQ)  2'd0;
     else if (link_down_reset_i)
       output_fifo_occupancy <= #(TCQ)  2'd0;
     else
       if ((in_data_valid_i & ~output_fifo_full) &
       ~((downstream_ready_i[3] | ~out_data_valid_o) &
         ~output_fifo_empty))
     output_fifo_occupancy <= #(TCQ) output_fifo_occupancy + 2'd1;
       else
     if (~(in_data_valid_i & ~output_fifo_full) &
         ((downstream_ready_i[3] | ~out_data_valid_o) &
          ~output_fifo_empty))
       output_fifo_occupancy <= #(TCQ) output_fifo_occupancy - 2'd1;
   
   assign output_fifo_full = output_fifo_occupancy[1];
   assign output_fifo_empty = (output_fifo_occupancy == 2'b00);

   // Write data into FIFO.
   always @(posedge clk_i)
     if (~reset_n_i)
       begin
          m_axis_rq_tdata_first_reg <= #(TCQ) {OUT_DATA_WIDTH{1'b0}};
          m_axis_rq_tdata_second_reg <= #(TCQ) {OUT_DATA_WIDTH{1'b0}};
          m_axis_rq_tkeep_first_reg <= #(TCQ) {TKEEP_WIDTH{1'b0}};
          m_axis_rq_tkeep_second_reg <= #(TCQ) {TKEEP_WIDTH{1'b0}};
          m_axis_rq_tuser_first_reg <= #(TCQ) {TUSER_WIDTH{1'b0}};
          m_axis_rq_tuser_second_reg <= #(TCQ) {TUSER_WIDTH{1'b0}};
          m_axis_rq_tlast_first_reg <= #(TCQ) 1'b0;
          m_axis_rq_tlast_second_reg <= #(TCQ) 1'b0;
       end
     else
        if (in_data_valid_i & ~output_fifo_full)
      begin
        case(output_fifo_write_ptr)
          1'b0:
         begin
            m_axis_rq_tdata_first_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH-1:0];
            m_axis_rq_tkeep_first_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH-1:OUT_DATA_WIDTH];
            m_axis_rq_tuser_first_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH+TUSER_WIDTH-1:OUT_DATA_WIDTH+TKEEP_WIDTH];
            m_axis_rq_tlast_first_reg <= #(TCQ) in_data_i[IN_DATA_WIDTH-1];
         end
           default:
         begin
            m_axis_rq_tdata_second_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH-1:0];
            m_axis_rq_tkeep_second_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH-1:OUT_DATA_WIDTH];
            m_axis_rq_tuser_second_reg <= #(TCQ) in_data_i[OUT_DATA_WIDTH+TKEEP_WIDTH+TUSER_WIDTH-1:OUT_DATA_WIDTH+TKEEP_WIDTH];
            m_axis_rq_tlast_second_reg <= #(TCQ) in_data_i[IN_DATA_WIDTH-1];
         end
         endcase // case(output_fifo_write_ptr)
        end // if (in_data_valid_i & ~output_fifo_full)
   
   // Output registers
   assign output_reg_mux_sel = output_fifo_read_ptr;

   always @(posedge clk_i)
     if (~reset_n_i)
       begin
      out_data_o <= #(TCQ)  {OUT_DATA_WIDTH{1'b0}};
      out_tuser_o <= #(TCQ)  {TUSER_WIDTH{1'b0}};
      out_tkeep_o <= #(TCQ)  {TKEEP_WIDTH{1'b0}};
      out_tlast_o <= #(TCQ)  1'b0;
       end
     else
       begin
      if (~out_data_valid_o | downstream_ready_i[0])
        begin
           case(output_reg_mux_sel)
         1'b0:
           begin
              out_data_o[127:0] <= #(TCQ)  m_axis_rq_tdata_first_reg[127:0];
           end
         default:
           begin
              out_data_o[127:0] <= #(TCQ)  m_axis_rq_tdata_second_reg[127:0];
           end
           endcase // case(output_reg_mux_sel)
        end // if (~out_data_valid_o | downstream_ready_i[0])

      if (~out_data_valid_o | downstream_ready_i[1])
        begin
           case(output_reg_mux_sel)
         1'b0:
           begin
              out_data_o[255:128] <= #(TCQ)  m_axis_rq_tdata_first_reg[255:128];
           end
         default:
           begin
              out_data_o[255:128] <= #(TCQ)  m_axis_rq_tdata_second_reg[255:128];
           end
           endcase // case(output_reg_mux_sel)
        end // if (~out_data_valid_o | downstream_ready_i[1])
      
      if (~out_data_valid_o | downstream_ready_i[2])
        begin
           case(output_reg_mux_sel)
         1'b0:
           begin
              out_tuser_o <= #(TCQ)  m_axis_rq_tuser_first_reg;
           end
         default:
           begin
              out_tuser_o <= #(TCQ)  m_axis_rq_tuser_second_reg;
           end
           endcase // case(output_reg_mux_sel)
        end // if (~out_data_valid_o | downstream_ready_i[2])
      
      if (~out_data_valid_o | downstream_ready_i[3])
        begin
           case(output_reg_mux_sel)
         1'b0:         
           begin
              out_tkeep_o <= #(TCQ)  m_axis_rq_tkeep_first_reg;
              out_tlast_o <= #(TCQ)  m_axis_rq_tlast_first_reg;
           end
         default:
           begin
              out_tkeep_o <= #(TCQ)  m_axis_rq_tkeep_second_reg;
              out_tlast_o <= #(TCQ)  m_axis_rq_tlast_second_reg;
           end
           endcase // case(output_reg_mux_sel)
        end // if (~out_data_valid_o | downstream_ready_i[3])
       end // else: !if(~reset_n_i)

   always @(posedge clk_i)
     if (~reset_n_i)
       out_data_valid_o <= #(TCQ) 1'b0;
     else
       if (~out_data_valid_o | downstream_ready_i[0])
     out_data_valid_o <= #(TCQ) ~output_fifo_empty;

endmodule // pcie_4_0_512b_rq_output_mux

//-----------------------------------------------------------------------------
//
// (c) Copyright 2012-2012 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//-----------------------------------------------------------------------------
//
// Project    : UltraScale+ FPGA PCI Express v4.0 Integrated Block
// File       : xp4_usp_smsw_512b_sync_fifo.v
// Version    : 1.1 
//-----------------------------------------------------------------------------
//--------------------------------------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)
module xp4_usp_smsw_512b_sync_fifo #
  (
   parameter TCQ = 100,
   parameter IMPL_TARGET = "SOFT",
   parameter AXISTEN_IF_EXT_512_INTFC_RAM_STYLE = "SRL",
   parameter FIFO_WIDTH = 512,
   parameter FIFO_DEPTH = 8,
   parameter FIFO_ALMOST_FULL_THRESHOLD = 5
   ) 
  (
    input  wire           clk_i // clock
   ,input  wire           reset_n_i // Reset
   ,input  wire           link_down_reset_i // Reset FIFO on link down

   ,input wire [FIFO_WIDTH-1:0] write_data_i
   ,input wire write_en_i
   ,input wire read_en_i
   ,output wire [FIFO_WIDTH-1:0] read_data_o
   ,output wire read_data_valid_o
   ,output reg fifo_almost_full
   );
   
   reg [2:0] write_ptr;
   reg [2:0] read_ptr;
   reg [3:0] fifo_occupancy;
   wire      fifo_empty;
   wire      fifo_full;

  integer    i;

   reg [FIFO_WIDTH-1:0] ram_array[FIFO_DEPTH-1:0];
   
  // SRL 16 should be inferred when RAM_STYLE = "SRL"
  generate 
    if (AXISTEN_IF_EXT_512_INTFC_RAM_STYLE =="SRL") 
      begin: srl_style_fifo

    // synthesis translate_off
    initial
          begin
        for (i=0; i < FIFO_DEPTH; i=i+1)
          ram_array[i] = 0;
      end
        // synthesis translate_on

  //Write to SRL inputs, and shift SRL
  always @(posedge clk_i)
      if (write_en_i & ~fifo_full)
        begin
      for (i= (FIFO_DEPTH-1); i>0; i=i-1)
        ram_array[i] <= #TCQ ram_array[i-1];
      ram_array[0]    <= #TCQ write_data_i;
        end

  //Maintain read pointer based on occupancy of the FIFO.
  // Read pointer points to the highest index of full locations.
   always @(posedge clk_i)
     if (~reset_n_i)
       read_ptr <= #TCQ 3'd0;
     else if (link_down_reset_i)
       read_ptr <= #TCQ 3'd0;
     else if (write_en_i && ~fifo_full &&
          (~(read_en_i & ~fifo_empty)))
       // Write but no read
       begin
     if (~fifo_empty)
       read_ptr <= #TCQ read_ptr + 3'd1;
       end
     else if ((~(write_en_i & ~fifo_full)) &&
          read_en_i && ~fifo_empty &&
          (read_ptr != 3'd0))
       // Read but no write
       read_ptr <= #TCQ read_ptr - 3'd1;

     assign    read_data_o = ram_array[read_ptr];
   end // block: srl_style_fifo
    else
      begin
   // Write pointer
   always @(posedge clk_i)
     if (~reset_n_i)
       write_ptr <= #TCQ 3'd0;
     else if (link_down_reset_i)
       write_ptr <= #TCQ 3'd0;
     else if (write_en_i & ~fifo_full)
       begin
      if (write_ptr == FIFO_DEPTH-1)
        write_ptr <= #TCQ 3'd0;
      else
        write_ptr <= #TCQ write_ptr + 3'd1;
       end
   always @(posedge clk_i)
     if (write_en_i & ~fifo_full)
       ram_array[write_ptr] <= #TCQ write_data_i;

   // Read pointer
   always @(posedge clk_i)
     if (~reset_n_i)
       read_ptr <= #TCQ 3'd0;
     else if (link_down_reset_i)
       read_ptr <= #TCQ 3'd0;
     else if (read_en_i & ~fifo_empty)
       begin
      if (read_ptr == FIFO_DEPTH-1)
        read_ptr <= #TCQ 3'd0;
      else
        read_ptr <= #TCQ read_ptr + 3'd1;
       end
    assign    read_data_o = ram_array[read_ptr];

    end // else: !if(AXISTEN_IF_EXT_512_INTFC_RAM_STYLE =="SRL")
  endgenerate

   // Maintain FIFO occupancy
   always @(posedge clk_i)
     if (~reset_n_i)
       fifo_occupancy <= #TCQ 4'd0;
     else if (link_down_reset_i)
       fifo_occupancy <= #TCQ 4'd0;
     else if (write_en_i & ~fifo_full &
          ~(read_en_i & ~fifo_empty))
       fifo_occupancy <= #TCQ fifo_occupancy + 4'd1;
     else if (~(write_en_i & ~fifo_full) &
          read_en_i & ~fifo_empty)
       fifo_occupancy <= #TCQ fifo_occupancy - 4'd1;

   always @(posedge clk_i)
     if (~reset_n_i)
       fifo_almost_full <= #TCQ 1'b0;
     else
       fifo_almost_full <= #TCQ (fifo_occupancy >= FIFO_ALMOST_FULL_THRESHOLD);

   assign    fifo_empty = (fifo_occupancy == 4'd0);
   assign    fifo_full = (fifo_occupancy == FIFO_DEPTH);
   assign    read_data_valid_o = ~fifo_empty;

endmodule // pcie_4_0_512b_sync_fifo

//
// Gen4 Specific Module - GEN4
//

