.GT_REFCLK0(gt_refclk0_out),

.apb3clk(iffctrlq0apb3clk),
.axisclk(iffctrlq0axisclk),

.apb3psel(iffctrlq0psel),
.apb3paddr(iffctrlq0paddr),
.apb3prdata(iffctrlq0prdata),
.apb3pready(iffctrlq0pready),
.apb3pwdata(iffctrlq0pwdata),
.apb3pwrite(iffctrlq0pwrite),
.apb3penable(iffctrlq0penable),
.apb3presetn(iffctrlq0presetn),
.apb3pslverr(iffctrlq0pslverr),

.bgpdb(iffctrlq0bgpwrdnb),
.bgbypassb(iffctrlq0bgbypass),
.bgrcalovrd(iffctrlq0bgrcalctl),
.bgmonitorenb(iffctrlq0bgtesten),
.bgrcalovrdenb(iffctrlq0bgrcalovrdenb),

.ch0_rxdata(iffcq00rxdata),
.ch0_rxrate(iffcq00rxrate),
.ch0_txdata(iffcq00txdata),
.ch0_txrate(iffcq00txrate),
.ch0_bufgtce(iffcq00bufgtce),
.ch0_gtrsvd(iffcq00pinrsrvd),
.ch0_pcierstb(iffcq00perstb),
.ch0_rxctrl0(iffcq00rxctrl0),
.ch0_rxctrl1(iffcq00rxctrl1),
.ch0_rxctrl2(iffcq00rxctrl2),
.ch0_rxctrl3(iffcq00rxctrl3),
.ch0_rxlpmen(iffcq00rxlpmen),
.ch0_rxpkdet(q0_ch0_rxpkdet),
.ch0_rxqpien(iffcq00rxqpien),
.ch0_rxslide(iffcq00rxslide),
.ch0_rxvalid(iffcq00rxvalid),
.ch0_tstclk0(iffcq00tstclk0),
.ch0_tstclk1(iffcq00tstclk1),
.ch0_txctrl0(iffcq00txctrl0),
.ch0_txctrl1(iffcq00txctrl1),
.ch0_txctrl2(iffcq00txctrl2),
.ch0_txpippmen(iffcq00enppm),
.ch0_txswing(iffcq00txswing),
.ch0_rxpd(iffcq00rxpowerdown),
.ch0_txpd(iffcq00txpowerdown),
.ch0_bufgtdiv(iffcq00bufgtdiv),
.ch0_bufgtrst(iffcq00bufgtrst),
.ch0_iloreset(iffcq00iloreset),
.ch0_loopback(iffcq00loopback),
.ch0_phyready(iffcq00phyready),
.ch0_rxcdrhold(iffcq00cdrhold),
.ch0_rxcdrlock(iffcq00cdrlock),
.ch0_rxheader(iffcq00rxheader),
.ch0_rxlatclk(iffcq00rxlatclk),
.ch0_rxoutclk(q0_ch0_rxoutclk),
.ch0_rxstatus(iffcq00rxstatus),
.ch0_rxusrclk(iffcq00rxusrclk),
.ch0_txcomsas(iffcq00txcomsas),
.ch0_txdeemph(iffcq00txdeemph),
.ch0_txheader(iffcq00txheader),
.ch0_txlatclk(iffcq00txlatclk),
.ch0_txmargin(iffcq00txmargin),
.ch0_txoutclk(q0_ch0_txoutclk),
.ch0_txusrclk(iffcq00txusrclk),
.ch0_dfehold(iffcq00aptexthold),
.ch0_rxuserrdy(iffcq00rxusrrdy),
.ch0_txuserrdy(iffcq00txusrrdy),
.ch0_cdrfreqos(iffcq00cdrfreqos),
.ch0_cdrstepsq(iffcq00cdrstepsq),
.ch0_cdrstepsx(iffcq00cdrstepsx),
.ch0_dfeovrd(iffcq00aptoverwren),
.ch0_dmonitorclk(iffcq00dmonclk),
.ch0_dmonitorout(iffcq00dmonout),
.ch0_gtrxreset(iffcq00gtrxreset),
.ch0_gttxreset(iffcq00gttxreset),
.ch0_pcsrsvdin(iffcq00pcsrsvdin),
.ch0_phystatus(iffcq00phystatus),
.ch0_rxchbondi(iffcq00rxchbondi),
.ch0_rxchbondo(iffcq00rxchbondo),
.ch0_rxprbserr(iffcq00rxprbserr),
.ch0_rxprbssel(iffcq00rxprbssel),
.ch0_rxqpisenn(iffcq00rxqpisenn),
.ch0_rxqpisenp(iffcq00rxqpisenp),
.ch0_txcominit(iffcq00txcominit),
.ch0_txcomwake(iffcq00txcomwake),
.ch0_txdccdone(iffcq00txdccdone),
.ch0_txdiffctrl(iffcq00txdrvamp),
.ch0_txinhibit(iffcq00txinhibit),
.ch0_txpisopd(iffcq00txserpwrdn),
.ch0_txprbssel(iffcq00txprbssel),
.ch0_txqpisenn(iffcq00txqpisenn),
.ch0_txqpisenp(iffcq00txqpisenp),
.ch0_clkrsvd0(iffcq00ckpinrsrvd0),
.ch0_clkrsvd1(iffcq00ckpinrsrvd1),
.ch0_pinrsvdas(iffcq00pinrsrvdas),
.ch0_rxcdrovrden(iffcq00cdrovren),
.ch0_rxosintdone(iffcq00cfokdone),
.ch0_txprecursor(iffcq00txemppre),
.ch0_cdrstepdir(iffcq00cdrstepdir),
.ch0_pcsrsvdout(iffcq00pcsrsvdout),
.ch0_refdebugout(iffcq00refclkpma),
.ch0_rxcdrreset(iffcq00cdrphreset),
.ch0_rxcommadet(iffcq00rxcommadet),
.ch0_rxcomsasdet(iffcq00comsasdet),
.ch0_rxelecidle(iffcq00rxelecidle),
.ch0_rxoobreset(iffcq00rxoobreset),
.ch0_rxpolarity(iffcq00rxpolarity),
.ch0_rxsliderdy(iffcq00rxsliderdy),
.ch0_rxslipdone(iffcq00rxslipdone),
.ch0_rxsyncdone(iffcq00rxsyncdone),
.ch0_txelecidle(iffcq00txelecidle),
.ch0_txpolarity(iffcq00txpolarity),
.ch0_txpostcursor(iffcq00txemppos),
.ch0_txsequence(iffcq00txsequence),
.ch0_txsyncdone(iffcq00txsyncdone),
.ch0_cdrbmcdrreq(iffcq00cdrbmcdreq),
.ch0_rxclkcorcnt(iffcq00rxckcorcnt),
.ch0_txmaincursor(iffcq00txempmain),
.ch0_bufgtcemask(iffcq00bufgtcemask),
.ch0_cdrincpctrl(iffcq00cdrincpctrl),
.ch0_rxbufstatus(iffcq00rxbufstatus),
.ch0_rxcdrphdone(iffcq00rxcdrphdone),
.ch0_rxcominitdet(iffcq00cominitdet),
.ch0_rxcomwakedet(iffcq00comwakedet),
.ch0_rxdapireset(iffcq00rxdapireset),
.ch0_rxdatavalid(iffcq00rxdatavalid),
.ch0_rxresetdone(iffcq00rxresetdone),
.ch0_rxresetmode(iffcq00rxresetmode),
.ch0_rxsyncallin(iffcq00rxsyncallin),
.ch0_txbufstatus(iffcq00txbufstatus),
.ch0_txcomfinish(iffcq00txcomfinish),
.ch0_txdapireset(iffcq00txdapireset),
.ch0_txoneszeros(iffcq00txoneszeros),
.ch0_txqpibiasen(iffcq00txqpibiasen),
.ch0_txqpiweakpu(iffcq00txqpiweakpu),
.ch0_txresetdone(iffcq00txresetdone),
.ch0_txresetmode(iffcq00txresetmode),
.ch0_txsyncallin(iffcq00txsyncallin),
.ch0_rxphdlypd(iffcq00rxphasealignpd),
.ch0_txphdlypd(iffcq00txphasealignpd),
.ch0_bufgtrstmask(iffcq00bufgtrstmask),
.ch0_eyescanreset(iffcq00eyescanreset),
.ch0_hsdppcsreset(iffcq00hsdppcsreset),
.ch0_iloresetdone(iffcq00iloresetdone),
.ch0_iloresetmask(iffcq00iloresetmask),
.ch0_rxdebugpcsout(iffcq00rxoutpcsclk),
.ch0_rxeqtraining(iffcq00rxeqtraining),
.ch0_rxphdlyreset(iffcq00rxphdlyreset),
.ch0_rxprbslocked(iffcq00rxprbslocked),
.ch0_rxstartofseq(iffcq00rxstartofseq),
.ch0_txdebugpcsout(iffcq00txoutpcsclk),
.ch0_txphdlyreset(iffcq00txphdlyreset),
.ch0_rxmstreset(iffctrlq0mstrxreset[0]),
.ch0_txmstreset(iffctrlq0msttxreset[0]),
.ch0_dmonfiforeset(iffcq00dmonfiforeset),
.ch0_rx10gstat(iffcq00rxethernetstatout),
.ch0_rxbyterealign(q0_ch0_rxbyterealign),
.ch0_rxchanbondseq(iffcq00rxchanbondseq),
.ch0_rxchanrealign(iffcq00rxchanrealign),
.ch0_rxgearboxslip(iffcq00rxgearboxslip),
.ch0_rxheadervalid(iffcq00rxheadervalid),
.ch0_rxmldchainreq(iffcq00rxmldchainreq),
.ch0_rxtermination(iffcq00rxtermination),
.ch0_txmldchainreq(iffcq00txmldchainreq),
.ch0_txpippmstepsize(iffcq00stepsizeppm),
.ch0_txswingoutlow(iffcq00txswingoutlow),
.ch0_rxphalignerr(iffcq00rxphasealignerr),
.ch0_rxphalignreq(iffcq00rxphasealignreq),
.ch0_txphalignerr(iffcq00txphasealignerr),
.ch0_txphalignreq(iffcq00txphasealignreq),
.ch0_txphdlytstclk(iffcq00tcoclkfsmfrout),
.ch0_dmonitoroutclk(q0_ch0_dmonitoroutclk),
.ch0_eyescantrigger(iffcq00eyescantrigger),
.ch0_resetexception(iffcq00resetexception),
.ch0_rxchanisaligned(iffcq00rxchisaligned),
.ch0_rxdlyalignerr(iffcq00rxdelayalignerr),
.ch0_rxdlyalignreq(iffcq00rxdelayalignreq),
.ch0_rxmldchaindone(iffcq00rxmldchaindone),
.ch0_rxpcsresetmask(iffcq00rxpcsresetmask),
.ch0_rxpmaresetdone(iffcq00rxpmaresetdone),
.ch0_rxpmaresetmask(iffcq00rxpmaresetmask),
.ch0_rxprbscntreset(iffcq00rxprbscntreset),
.ch0_rxprogdivreset(iffcq00rxprogdivreset),
.ch0_txdetectrx(iffcq00txdetectrxloopback),
.ch0_txdlyalignerr(iffcq00txdelayalignerr),
.ch0_txdlyalignreq(iffcq00txdelayalignreq),
.ch0_txmldchaindone(iffcq00txmldchaindone),
.ch0_txpcsresetmask(iffcq00txpcsresetmask),
.ch0_txpicodereset(iffcq00txtxpicodereset),
.ch0_txpmaresetdone(iffcq00txpmaresetdone),
.ch0_txpmaresetmask(iffcq00txpmaresetmask),
.ch0_txprbsforceerr(iffcq00txprbsforceerr),
.ch0_txprogdivreset(iffcq00txprogdivreset),
.ch0_txswingouthigh(iffcq00txswingouthigh),
.ch0_rxphaligndone(iffcq00rxphasealigndone),
.ch0_txphaligndone(iffcq00txphasealigndone),
.ch0_rxbyteisaligned(iffcq00rxbyteisaligned),
.ch0_rxdapicodereset(iffcq00rxdapicodereset),
.ch0_rxdapiresetdone(iffcq00rxdapiresetdone),
.ch0_rxdapiresetmask(iffcq00rxdapiresetmask),
.ch0_rxfinealigndone(iffcq00rxfinealigndone),
.ch0_rxphshift180(iffcq00rxphaseshift180req),
.ch0_txdapicodereset(iffcq00txdapicodereset),
.ch0_txdapiresetdone(iffcq00txdapiresetdone),
.ch0_txdapiresetmask(iffcq00txdapiresetmask),
.ch0_txphalignoutrsvd(iffcq00txchicooutrsvd),
.ch0_txphshift180(iffcq00txphaseshift180req),
.ch0_txpicodeovrden(iffcq00txtxpicodeovrden),
.ch0_rxphsetinitreq(iffcq00rxphasesetinitreq),
.ch0_txphsetinitreq(iffcq00txphasesetinitreq),
.ch0_eyescandataerror(iffcq00eyescandataerror),
.ch0_rxdapicodeovrden(iffcq00rxdapicodeovrden),
.ch0_rxmlfinealignreq(iffcq00rxmlfinealignreq),
.ch0_txdapicodeovrden(iffcq00txdapicodeovrden),
.ch0_rxmstresetdone(iffctrlq0mstrxresetdone[0]),
.ch0_rxphsetinitdone(iffcq00rxphasesetinitdone),
.ch0_txmstresetdone(iffctrlq0msttxresetdone[0]),
.ch0_txphsetinitdone(iffcq00txphasesetinitdone),
.ch0_rxdlyalignprog(iffcq00rxdelayalignprogress),
.ch0_rxphalignresetmask(iffcq00rxchicoresetmask),
.ch0_txdlyalignprog(iffcq00txdelayalignprogress),
.ch0_txpausedelayalign(iffcq00txpausedelayalign),
.ch0_txphalignresetmask(iffcq00txchicoresetmask),
.ch0_xpipe5_pipeline_en(iffcq00xpipe5pipelineen),
.ch0_phyesmadaptsave(iffcq00phyesmadaptationsave),
.ch0_rxphshift180done(iffcq00rxphaseshift180done),
.ch0_tx10gstat(iffcq00txethernetstattxlocalfault),
.ch0_txphshift180done(iffcq00txphaseshift180done),
.ch0_rxprogdivresetdone(iffcq00rxprogdivresetdone),
.ch0_rxsimplexphystatus(iffcq00rxsimplexphystatus),
.ch0_txprogdivresetdone(iffcq00txprogdivresetdone),
.ch0_txsimplexphystatus(iffcq00txsimplexphystatus),
.ch0_rxphdlyresetdone(iffcq00rxphasedelayresetdone),
.ch0_txphdlyresetdone(iffcq00txphasedelayresetdone),

.ch1_rxdata(iffcq01rxdata),
.ch1_rxrate(iffcq01rxrate),
.ch1_txdata(iffcq01txdata),
.ch1_txrate(iffcq01txrate),
.ch1_bufgtce(iffcq01bufgtce),
.ch1_gtrsvd(iffcq01pinrsrvd),
.ch1_pcierstb(iffcq01perstb),
.ch1_rxctrl0(iffcq01rxctrl0),
.ch1_rxctrl1(iffcq01rxctrl1),
.ch1_rxctrl2(iffcq01rxctrl2),
.ch1_rxctrl3(iffcq01rxctrl3),
.ch1_rxlpmen(iffcq01rxlpmen),
.ch1_rxpkdet(q0_ch1_rxpkdet),
.ch1_rxqpien(iffcq01rxqpien),
.ch1_rxslide(iffcq01rxslide),
.ch1_rxvalid(iffcq01rxvalid),
.ch1_tstclk0(iffcq01tstclk0),
.ch1_tstclk1(iffcq01tstclk1),
.ch1_txctrl0(iffcq01txctrl0),
.ch1_txctrl1(iffcq01txctrl1),
.ch1_txctrl2(iffcq01txctrl2),
.ch1_txpippmen(iffcq01enppm),
.ch1_txswing(iffcq01txswing),
.ch1_rxpd(iffcq01rxpowerdown),
.ch1_txpd(iffcq01txpowerdown),
.ch1_bufgtdiv(iffcq01bufgtdiv),
.ch1_bufgtrst(iffcq01bufgtrst),
.ch1_iloreset(iffcq01iloreset),
.ch1_loopback(iffcq01loopback),
.ch1_phyready(iffcq01phyready),
.ch1_rxcdrhold(iffcq01cdrhold),
.ch1_rxcdrlock(iffcq01cdrlock),
.ch1_rxheader(iffcq01rxheader),
.ch1_rxlatclk(iffcq01rxlatclk),
.ch1_rxoutclk(q0_ch1_rxoutclk),
.ch1_rxstatus(iffcq01rxstatus),
.ch1_rxusrclk(iffcq01rxusrclk),
.ch1_txcomsas(iffcq01txcomsas),
.ch1_txdeemph(iffcq01txdeemph),
.ch1_txheader(iffcq01txheader),
.ch1_txlatclk(iffcq01txlatclk),
.ch1_txmargin(iffcq01txmargin),
.ch1_txoutclk(q0_ch1_txoutclk),
.ch1_txusrclk(iffcq01txusrclk),
.ch1_dfehold(iffcq01aptexthold),
.ch1_rxuserrdy(iffcq01rxusrrdy),
.ch1_txuserrdy(iffcq01txusrrdy),
.ch1_cdrfreqos(iffcq01cdrfreqos),
.ch1_cdrstepsq(iffcq01cdrstepsq),
.ch1_cdrstepsx(iffcq01cdrstepsx),
.ch1_dfeovrd(iffcq01aptoverwren),
.ch1_dmonitorclk(iffcq01dmonclk),
.ch1_dmonitorout(iffcq01dmonout),
.ch1_gtrxreset(iffcq01gtrxreset),
.ch1_gttxreset(iffcq01gttxreset),
.ch1_pcsrsvdin(iffcq01pcsrsvdin),
.ch1_phystatus(iffcq01phystatus),
.ch1_rxchbondi(iffcq01rxchbondi),
.ch1_rxchbondo(iffcq01rxchbondo),
.ch1_rxprbserr(iffcq01rxprbserr),
.ch1_rxprbssel(iffcq01rxprbssel),
.ch1_rxqpisenn(iffcq01rxqpisenn),
.ch1_rxqpisenp(iffcq01rxqpisenp),
.ch1_txcominit(iffcq01txcominit),
.ch1_txcomwake(iffcq01txcomwake),
.ch1_txdccdone(iffcq01txdccdone),
.ch1_txdiffctrl(iffcq01txdrvamp),
.ch1_txinhibit(iffcq01txinhibit),
.ch1_txpisopd(iffcq01txserpwrdn),
.ch1_txprbssel(iffcq01txprbssel),
.ch1_txqpisenn(iffcq01txqpisenn),
.ch1_txqpisenp(iffcq01txqpisenp),
.ch1_clkrsvd0(iffcq01ckpinrsrvd0),
.ch1_clkrsvd1(iffcq01ckpinrsrvd1),
.ch1_pinrsvdas(iffcq01pinrsrvdas),
.ch1_rxcdrovrden(iffcq01cdrovren),
.ch1_rxosintdone(iffcq01cfokdone),
.ch1_txprecursor(iffcq01txemppre),
.ch1_cdrstepdir(iffcq01cdrstepdir),
.ch1_pcsrsvdout(iffcq01pcsrsvdout),
.ch1_refdebugout(iffcq01refclkpma),
.ch1_rxcdrreset(iffcq01cdrphreset),
.ch1_rxcommadet(iffcq01rxcommadet),
.ch1_rxcomsasdet(iffcq01comsasdet),
.ch1_rxelecidle(iffcq01rxelecidle),
.ch1_rxoobreset(iffcq01rxoobreset),
.ch1_rxpolarity(iffcq01rxpolarity),
.ch1_rxsliderdy(iffcq01rxsliderdy),
.ch1_rxslipdone(iffcq01rxslipdone),
.ch1_rxsyncdone(iffcq01rxsyncdone),
.ch1_txelecidle(iffcq01txelecidle),
.ch1_txpolarity(iffcq01txpolarity),
.ch1_txpostcursor(iffcq01txemppos),
.ch1_txsequence(iffcq01txsequence),
.ch1_txsyncdone(iffcq01txsyncdone),
.ch1_cdrbmcdrreq(iffcq01cdrbmcdreq),
.ch1_rxclkcorcnt(iffcq01rxckcorcnt),
.ch1_txmaincursor(iffcq01txempmain),
.ch1_bufgtcemask(iffcq01bufgtcemask),
.ch1_cdrincpctrl(iffcq01cdrincpctrl),
.ch1_rxbufstatus(iffcq01rxbufstatus),
.ch1_rxcdrphdone(iffcq01rxcdrphdone),
.ch1_rxcominitdet(iffcq01cominitdet),
.ch1_rxcomwakedet(iffcq01comwakedet),
.ch1_rxdapireset(iffcq01rxdapireset),
.ch1_rxdatavalid(iffcq01rxdatavalid),
.ch1_rxresetdone(iffcq01rxresetdone),
.ch1_rxresetmode(iffcq01rxresetmode),
.ch1_rxsyncallin(iffcq01rxsyncallin),
.ch1_txbufstatus(iffcq01txbufstatus),
.ch1_txcomfinish(iffcq01txcomfinish),
.ch1_txdapireset(iffcq01txdapireset),
.ch1_txoneszeros(iffcq01txoneszeros),
.ch1_txqpibiasen(iffcq01txqpibiasen),
.ch1_txqpiweakpu(iffcq01txqpiweakpu),
.ch1_txresetdone(iffcq01txresetdone),
.ch1_txresetmode(iffcq01txresetmode),
.ch1_txsyncallin(iffcq01txsyncallin),
.ch1_rxphdlypd(iffcq01rxphasealignpd),
.ch1_txphdlypd(iffcq01txphasealignpd),
.ch1_bufgtrstmask(iffcq01bufgtrstmask),
.ch1_eyescanreset(iffcq01eyescanreset),
.ch1_hsdppcsreset(iffcq01hsdppcsreset),
.ch1_iloresetdone(iffcq01iloresetdone),
.ch1_iloresetmask(iffcq01iloresetmask),
.ch1_rxdebugpcsout(iffcq01rxoutpcsclk),
.ch1_rxeqtraining(iffcq01rxeqtraining),
.ch1_rxphdlyreset(iffcq01rxphdlyreset),
.ch1_rxprbslocked(iffcq01rxprbslocked),
.ch1_rxstartofseq(iffcq01rxstartofseq),
.ch1_txdebugpcsout(iffcq01txoutpcsclk),
.ch1_txphdlyreset(iffcq01txphdlyreset),
.ch1_rxmstreset(iffctrlq0mstrxreset[1]),
.ch1_txmstreset(iffctrlq0msttxreset[1]),
.ch1_dmonfiforeset(iffcq01dmonfiforeset),
.ch1_rx10gstat(iffcq01rxethernetstatout),
.ch1_rxbyterealign(q0_ch1_rxbyterealign),
.ch1_rxchanbondseq(iffcq01rxchanbondseq),
.ch1_rxchanrealign(iffcq01rxchanrealign),
.ch1_rxgearboxslip(iffcq01rxgearboxslip),
.ch1_rxheadervalid(iffcq01rxheadervalid),
.ch1_rxmldchainreq(iffcq01rxmldchainreq),
.ch1_rxtermination(iffcq01rxtermination),
.ch1_txmldchainreq(iffcq01txmldchainreq),
.ch1_txpippmstepsize(iffcq01stepsizeppm),
.ch1_txswingoutlow(iffcq01txswingoutlow),
.ch1_rxphalignerr(iffcq01rxphasealignerr),
.ch1_rxphalignreq(iffcq01rxphasealignreq),
.ch1_txphalignerr(iffcq01txphasealignerr),
.ch1_txphalignreq(iffcq01txphasealignreq),
.ch1_txphdlytstclk(iffcq01tcoclkfsmfrout),
.ch1_dmonitoroutclk(q0_ch1_dmonitoroutclk),
.ch1_eyescantrigger(iffcq01eyescantrigger),
.ch1_resetexception(iffcq01resetexception),
.ch1_rxchanisaligned(iffcq01rxchisaligned),
.ch1_rxdlyalignerr(iffcq01rxdelayalignerr),
.ch1_rxdlyalignreq(iffcq01rxdelayalignreq),
.ch1_rxmldchaindone(iffcq01rxmldchaindone),
.ch1_rxpcsresetmask(iffcq01rxpcsresetmask),
.ch1_rxpmaresetdone(iffcq01rxpmaresetdone),
.ch1_rxpmaresetmask(iffcq01rxpmaresetmask),
.ch1_rxprbscntreset(iffcq01rxprbscntreset),
.ch1_rxprogdivreset(iffcq01rxprogdivreset),
.ch1_txdetectrx(iffcq01txdetectrxloopback),
.ch1_txdlyalignerr(iffcq01txdelayalignerr),
.ch1_txdlyalignreq(iffcq01txdelayalignreq),
.ch1_txmldchaindone(iffcq01txmldchaindone),
.ch1_txpcsresetmask(iffcq01txpcsresetmask),
.ch1_txpicodereset(iffcq01txtxpicodereset),
.ch1_txpmaresetdone(iffcq01txpmaresetdone),
.ch1_txpmaresetmask(iffcq01txpmaresetmask),
.ch1_txprbsforceerr(iffcq01txprbsforceerr),
.ch1_txprogdivreset(iffcq01txprogdivreset),
.ch1_txswingouthigh(iffcq01txswingouthigh),
.ch1_rxphaligndone(iffcq01rxphasealigndone),
.ch1_txphaligndone(iffcq01txphasealigndone),
.ch1_rxbyteisaligned(iffcq01rxbyteisaligned),
.ch1_rxdapicodereset(iffcq01rxdapicodereset),
.ch1_rxdapiresetdone(iffcq01rxdapiresetdone),
.ch1_rxdapiresetmask(iffcq01rxdapiresetmask),
.ch1_rxfinealigndone(iffcq01rxfinealigndone),
.ch1_rxphshift180(iffcq01rxphaseshift180req),
.ch1_txdapicodereset(iffcq01txdapicodereset),
.ch1_txdapiresetdone(iffcq01txdapiresetdone),
.ch1_txdapiresetmask(iffcq01txdapiresetmask),
.ch1_txphalignoutrsvd(iffcq01txchicooutrsvd),
.ch1_txphshift180(iffcq01txphaseshift180req),
.ch1_txpicodeovrden(iffcq01txtxpicodeovrden),
.ch1_rxphsetinitreq(iffcq01rxphasesetinitreq),
.ch1_txphsetinitreq(iffcq01txphasesetinitreq),
.ch1_eyescandataerror(iffcq01eyescandataerror),
.ch1_rxdapicodeovrden(iffcq01rxdapicodeovrden),
.ch1_rxmlfinealignreq(iffcq01rxmlfinealignreq),
.ch1_txdapicodeovrden(iffcq01txdapicodeovrden),
.ch1_rxmstresetdone(iffctrlq0mstrxresetdone[1]),
.ch1_rxphsetinitdone(iffcq01rxphasesetinitdone),
.ch1_txmstresetdone(iffctrlq0msttxresetdone[1]),
.ch1_txphsetinitdone(iffcq01txphasesetinitdone),
.ch1_rxdlyalignprog(iffcq01rxdelayalignprogress),
.ch1_rxphalignresetmask(iffcq01rxchicoresetmask),
.ch1_txdlyalignprog(iffcq01txdelayalignprogress),
.ch1_txpausedelayalign(iffcq01txpausedelayalign),
.ch1_txphalignresetmask(iffcq01txchicoresetmask),
.ch1_xpipe5_pipeline_en(iffcq01xpipe5pipelineen),
.ch1_phyesmadaptsave(iffcq01phyesmadaptationsave),
.ch1_rxphshift180done(iffcq01rxphaseshift180done),
.ch1_tx10gstat(iffcq01txethernetstattxlocalfault),
.ch1_txphshift180done(iffcq01txphaseshift180done),
.ch1_rxprogdivresetdone(iffcq01rxprogdivresetdone),
.ch1_rxsimplexphystatus(iffcq01rxsimplexphystatus),
.ch1_txprogdivresetdone(iffcq01txprogdivresetdone),
.ch1_txsimplexphystatus(iffcq01txsimplexphystatus),
.ch1_rxphdlyresetdone(iffcq01rxphasedelayresetdone),
.ch1_txphdlyresetdone(iffcq01txphasedelayresetdone),

.ch2_rxdata(iffcq02rxdata),
.ch2_rxrate(iffcq02rxrate),
.ch2_txdata(iffcq02txdata),
.ch2_txrate(iffcq02txrate),
.ch2_bufgtce(iffcq02bufgtce),
.ch2_gtrsvd(iffcq02pinrsrvd),
.ch2_pcierstb(iffcq02perstb),
.ch2_rxctrl0(iffcq02rxctrl0),
.ch2_rxctrl1(iffcq02rxctrl1),
.ch2_rxctrl2(iffcq02rxctrl2),
.ch2_rxctrl3(iffcq02rxctrl3),
.ch2_rxlpmen(iffcq02rxlpmen),
.ch2_rxpkdet(q0_ch2_rxpkdet),
.ch2_rxqpien(iffcq02rxqpien),
.ch2_rxslide(iffcq02rxslide),
.ch2_rxvalid(iffcq02rxvalid),
.ch2_tstclk0(iffcq02tstclk0),
.ch2_tstclk1(iffcq02tstclk1),
.ch2_txctrl0(iffcq02txctrl0),
.ch2_txctrl1(iffcq02txctrl1),
.ch2_txctrl2(iffcq02txctrl2),
.ch2_txpippmen(iffcq02enppm),
.ch2_txswing(iffcq02txswing),
.ch2_rxpd(iffcq02rxpowerdown),
.ch2_txpd(iffcq02txpowerdown),
.ch2_bufgtdiv(iffcq02bufgtdiv),
.ch2_bufgtrst(iffcq02bufgtrst),
.ch2_iloreset(iffcq02iloreset),
.ch2_loopback(iffcq02loopback),
.ch2_phyready(iffcq02phyready),
.ch2_rxcdrhold(iffcq02cdrhold),
.ch2_rxcdrlock(iffcq02cdrlock),
.ch2_rxheader(iffcq02rxheader),
.ch2_rxlatclk(iffcq02rxlatclk),
.ch2_rxoutclk(q0_ch2_rxoutclk),
.ch2_rxstatus(iffcq02rxstatus),
.ch2_rxusrclk(iffcq02rxusrclk),
.ch2_txcomsas(iffcq02txcomsas),
.ch2_txdeemph(iffcq02txdeemph),
.ch2_txheader(iffcq02txheader),
.ch2_txlatclk(iffcq02txlatclk),
.ch2_txmargin(iffcq02txmargin),
.ch2_txoutclk(q0_ch2_txoutclk),
.ch2_txusrclk(iffcq02txusrclk),
.ch2_dfehold(iffcq02aptexthold),
.ch2_rxuserrdy(iffcq02rxusrrdy),
.ch2_txuserrdy(iffcq02txusrrdy),
.ch2_cdrfreqos(iffcq02cdrfreqos),
.ch2_cdrstepsq(iffcq02cdrstepsq),
.ch2_cdrstepsx(iffcq02cdrstepsx),
.ch2_dfeovrd(iffcq02aptoverwren),
.ch2_dmonitorclk(iffcq02dmonclk),
.ch2_dmonitorout(iffcq02dmonout),
.ch2_gtrxreset(iffcq02gtrxreset),
.ch2_gttxreset(iffcq02gttxreset),
.ch2_pcsrsvdin(iffcq02pcsrsvdin),
.ch2_phystatus(iffcq02phystatus),
.ch2_rxchbondi(iffcq02rxchbondi),
.ch2_rxchbondo(iffcq02rxchbondo),
.ch2_rxprbserr(iffcq02rxprbserr),
.ch2_rxprbssel(iffcq02rxprbssel),
.ch2_rxqpisenn(iffcq02rxqpisenn),
.ch2_rxqpisenp(iffcq02rxqpisenp),
.ch2_txcominit(iffcq02txcominit),
.ch2_txcomwake(iffcq02txcomwake),
.ch2_txdccdone(iffcq02txdccdone),
.ch2_txdiffctrl(iffcq02txdrvamp),
.ch2_txinhibit(iffcq02txinhibit),
.ch2_txpisopd(iffcq02txserpwrdn),
.ch2_txprbssel(iffcq02txprbssel),
.ch2_txqpisenn(iffcq02txqpisenn),
.ch2_txqpisenp(iffcq02txqpisenp),
.ch2_clkrsvd0(iffcq02ckpinrsrvd0),
.ch2_clkrsvd1(iffcq02ckpinrsrvd1),
.ch2_pinrsvdas(iffcq02pinrsrvdas),
.ch2_rxcdrovrden(iffcq02cdrovren),
.ch2_rxosintdone(iffcq02cfokdone),
.ch2_txprecursor(iffcq02txemppre),
.ch2_cdrstepdir(iffcq02cdrstepdir),
.ch2_pcsrsvdout(iffcq02pcsrsvdout),
.ch2_refdebugout(iffcq02refclkpma),
.ch2_rxcdrreset(iffcq02cdrphreset),
.ch2_rxcommadet(iffcq02rxcommadet),
.ch2_rxcomsasdet(iffcq02comsasdet),
.ch2_rxelecidle(iffcq02rxelecidle),
.ch2_rxoobreset(iffcq02rxoobreset),
.ch2_rxpolarity(iffcq02rxpolarity),
.ch2_rxsliderdy(iffcq02rxsliderdy),
.ch2_rxslipdone(iffcq02rxslipdone),
.ch2_rxsyncdone(iffcq02rxsyncdone),
.ch2_txelecidle(iffcq02txelecidle),
.ch2_txpolarity(iffcq02txpolarity),
.ch2_txpostcursor(iffcq02txemppos),
.ch2_txsequence(iffcq02txsequence),
.ch2_txsyncdone(iffcq02txsyncdone),
.ch2_cdrbmcdrreq(iffcq02cdrbmcdreq),
.ch2_rxclkcorcnt(iffcq02rxckcorcnt),
.ch2_txmaincursor(iffcq02txempmain),
.ch2_bufgtcemask(iffcq02bufgtcemask),
.ch2_cdrincpctrl(iffcq02cdrincpctrl),
.ch2_rxbufstatus(iffcq02rxbufstatus),
.ch2_rxcdrphdone(iffcq02rxcdrphdone),
.ch2_rxcominitdet(iffcq02cominitdet),
.ch2_rxcomwakedet(iffcq02comwakedet),
.ch2_rxdapireset(iffcq02rxdapireset),
.ch2_rxdatavalid(iffcq02rxdatavalid),
.ch2_rxresetdone(iffcq02rxresetdone),
.ch2_rxresetmode(iffcq02rxresetmode),
.ch2_rxsyncallin(iffcq02rxsyncallin),
.ch2_txbufstatus(iffcq02txbufstatus),
.ch2_txcomfinish(iffcq02txcomfinish),
.ch2_txdapireset(iffcq02txdapireset),
.ch2_txoneszeros(iffcq02txoneszeros),
.ch2_txqpibiasen(iffcq02txqpibiasen),
.ch2_txqpiweakpu(iffcq02txqpiweakpu),
.ch2_txresetdone(iffcq02txresetdone),
.ch2_txresetmode(iffcq02txresetmode),
.ch2_txsyncallin(iffcq02txsyncallin),
.ch2_rxphdlypd(iffcq02rxphasealignpd),
.ch2_txphdlypd(iffcq02txphasealignpd),
.ch2_bufgtrstmask(iffcq02bufgtrstmask),
.ch2_eyescanreset(iffcq02eyescanreset),
.ch2_hsdppcsreset(iffcq02hsdppcsreset),
.ch2_iloresetdone(iffcq02iloresetdone),
.ch2_iloresetmask(iffcq02iloresetmask),
.ch2_rxdebugpcsout(iffcq02rxoutpcsclk),
.ch2_rxeqtraining(iffcq02rxeqtraining),
.ch2_rxphdlyreset(iffcq02rxphdlyreset),
.ch2_rxprbslocked(iffcq02rxprbslocked),
.ch2_rxstartofseq(iffcq02rxstartofseq),
.ch2_txdebugpcsout(iffcq02txoutpcsclk),
.ch2_txphdlyreset(iffcq02txphdlyreset),
.ch2_rxmstreset(iffctrlq0mstrxreset[2]),
.ch2_txmstreset(iffctrlq0msttxreset[2]),
.ch2_dmonfiforeset(iffcq02dmonfiforeset),
.ch2_rx10gstat(iffcq02rxethernetstatout),
.ch2_rxbyterealign(q0_ch2_rxbyterealign),
.ch2_rxchanbondseq(iffcq02rxchanbondseq),
.ch2_rxchanrealign(iffcq02rxchanrealign),
.ch2_rxgearboxslip(iffcq02rxgearboxslip),
.ch2_rxheadervalid(iffcq02rxheadervalid),
.ch2_rxmldchainreq(iffcq02rxmldchainreq),
.ch2_rxtermination(iffcq02rxtermination),
.ch2_txmldchainreq(iffcq02txmldchainreq),
.ch2_txpippmstepsize(iffcq02stepsizeppm),
.ch2_txswingoutlow(iffcq02txswingoutlow),
.ch2_rxphalignerr(iffcq02rxphasealignerr),
.ch2_rxphalignreq(iffcq02rxphasealignreq),
.ch2_txphalignerr(iffcq02txphasealignerr),
.ch2_txphalignreq(iffcq02txphasealignreq),
.ch2_txphdlytstclk(iffcq02tcoclkfsmfrout),
.ch2_dmonitoroutclk(q0_ch2_dmonitoroutclk),
.ch2_eyescantrigger(iffcq02eyescantrigger),
.ch2_resetexception(iffcq02resetexception),
.ch2_rxchanisaligned(iffcq02rxchisaligned),
.ch2_rxdlyalignerr(iffcq02rxdelayalignerr),
.ch2_rxdlyalignreq(iffcq02rxdelayalignreq),
.ch2_rxmldchaindone(iffcq02rxmldchaindone),
.ch2_rxpcsresetmask(iffcq02rxpcsresetmask),
.ch2_rxpmaresetdone(iffcq02rxpmaresetdone),
.ch2_rxpmaresetmask(iffcq02rxpmaresetmask),
.ch2_rxprbscntreset(iffcq02rxprbscntreset),
.ch2_rxprogdivreset(iffcq02rxprogdivreset),
.ch2_txdetectrx(iffcq02txdetectrxloopback),
.ch2_txdlyalignerr(iffcq02txdelayalignerr),
.ch2_txdlyalignreq(iffcq02txdelayalignreq),
.ch2_txmldchaindone(iffcq02txmldchaindone),
.ch2_txpcsresetmask(iffcq02txpcsresetmask),
.ch2_txpicodereset(iffcq02txtxpicodereset),
.ch2_txpmaresetdone(iffcq02txpmaresetdone),
.ch2_txpmaresetmask(iffcq02txpmaresetmask),
.ch2_txprbsforceerr(iffcq02txprbsforceerr),
.ch2_txprogdivreset(iffcq02txprogdivreset),
.ch2_txswingouthigh(iffcq02txswingouthigh),
.ch2_rxphaligndone(iffcq02rxphasealigndone),
.ch2_txphaligndone(iffcq02txphasealigndone),
.ch2_rxbyteisaligned(iffcq02rxbyteisaligned),
.ch2_rxdapicodereset(iffcq02rxdapicodereset),
.ch2_rxdapiresetdone(iffcq02rxdapiresetdone),
.ch2_rxdapiresetmask(iffcq02rxdapiresetmask),
.ch2_rxfinealigndone(iffcq02rxfinealigndone),
.ch2_rxphshift180(iffcq02rxphaseshift180req),
.ch2_txdapicodereset(iffcq02txdapicodereset),
.ch2_txdapiresetdone(iffcq02txdapiresetdone),
.ch2_txdapiresetmask(iffcq02txdapiresetmask),
.ch2_txphalignoutrsvd(iffcq02txchicooutrsvd),
.ch2_txphshift180(iffcq02txphaseshift180req),
.ch2_txpicodeovrden(iffcq02txtxpicodeovrden),
.ch2_rxphsetinitreq(iffcq02rxphasesetinitreq),
.ch2_txphsetinitreq(iffcq02txphasesetinitreq),
.ch2_eyescandataerror(iffcq02eyescandataerror),
.ch2_rxdapicodeovrden(iffcq02rxdapicodeovrden),
.ch2_rxmlfinealignreq(iffcq02rxmlfinealignreq),
.ch2_txdapicodeovrden(iffcq02txdapicodeovrden),
.ch2_rxmstresetdone(iffctrlq0mstrxresetdone[2]),
.ch2_rxphsetinitdone(iffcq02rxphasesetinitdone),
.ch2_txmstresetdone(iffctrlq0msttxresetdone[2]),
.ch2_txphsetinitdone(iffcq02txphasesetinitdone),
.ch2_rxdlyalignprog(iffcq02rxdelayalignprogress),
.ch2_rxphalignresetmask(iffcq02rxchicoresetmask),
.ch2_txdlyalignprog(iffcq02txdelayalignprogress),
.ch2_txpausedelayalign(iffcq02txpausedelayalign),
.ch2_txphalignresetmask(iffcq02txchicoresetmask),
.ch2_xpipe5_pipeline_en(iffcq02xpipe5pipelineen),
.ch2_phyesmadaptsave(iffcq02phyesmadaptationsave),
.ch2_rxphshift180done(iffcq02rxphaseshift180done),
.ch2_tx10gstat(iffcq02txethernetstattxlocalfault),
.ch2_txphshift180done(iffcq02txphaseshift180done),
.ch2_rxprogdivresetdone(iffcq02rxprogdivresetdone),
.ch2_rxsimplexphystatus(iffcq02rxsimplexphystatus),
.ch2_txprogdivresetdone(iffcq02txprogdivresetdone),
.ch2_txsimplexphystatus(iffcq02txsimplexphystatus),
.ch2_rxphdlyresetdone(iffcq02rxphasedelayresetdone),
.ch2_txphdlyresetdone(iffcq02txphasedelayresetdone),

.ch3_rxdata(iffcq03rxdata),
.ch3_rxrate(iffcq03rxrate),
.ch3_txdata(iffcq03txdata),
.ch3_txrate(iffcq03txrate),
.ch3_bufgtce(iffcq03bufgtce),
.ch3_gtrsvd(iffcq03pinrsrvd),
.ch3_pcierstb(iffcq03perstb),
.ch3_rxctrl0(iffcq03rxctrl0),
.ch3_rxctrl1(iffcq03rxctrl1),
.ch3_rxctrl2(iffcq03rxctrl2),
.ch3_rxctrl3(iffcq03rxctrl3),
.ch3_rxlpmen(iffcq03rxlpmen),
.ch3_rxpkdet(q0_ch3_rxpkdet),
.ch3_rxqpien(iffcq03rxqpien),
.ch3_rxslide(iffcq03rxslide),
.ch3_rxvalid(iffcq03rxvalid),
.ch3_tstclk0(iffcq03tstclk0),
.ch3_tstclk1(iffcq03tstclk1),
.ch3_txctrl0(iffcq03txctrl0),
.ch3_txctrl1(iffcq03txctrl1),
.ch3_txctrl2(iffcq03txctrl2),
.ch3_txpippmen(iffcq03enppm),
.ch3_txswing(iffcq03txswing),
.ch3_rxpd(iffcq03rxpowerdown),
.ch3_txpd(iffcq03txpowerdown),
.ch3_bufgtdiv(iffcq03bufgtdiv),
.ch3_bufgtrst(iffcq03bufgtrst),
.ch3_iloreset(iffcq03iloreset),
.ch3_loopback(iffcq03loopback),
.ch3_phyready(iffcq03phyready),
.ch3_rxcdrhold(iffcq03cdrhold),
.ch3_rxcdrlock(iffcq03cdrlock),
.ch3_rxheader(iffcq03rxheader),
.ch3_rxlatclk(iffcq03rxlatclk),
.ch3_rxoutclk(q0_ch3_rxoutclk),
.ch3_rxstatus(iffcq03rxstatus),
.ch3_rxusrclk(iffcq03rxusrclk),
.ch3_txcomsas(iffcq03txcomsas),
.ch3_txdeemph(iffcq03txdeemph),
.ch3_txheader(iffcq03txheader),
.ch3_txlatclk(iffcq03txlatclk),
.ch3_txmargin(iffcq03txmargin),
.ch3_txoutclk(q0_ch3_txoutclk),
.ch3_txusrclk(iffcq03txusrclk),
.ch3_dfehold(iffcq03aptexthold),
.ch3_rxuserrdy(iffcq03rxusrrdy),
.ch3_txuserrdy(iffcq03txusrrdy),
.ch3_cdrfreqos(iffcq03cdrfreqos),
.ch3_cdrstepsq(iffcq03cdrstepsq),
.ch3_cdrstepsx(iffcq03cdrstepsx),
.ch3_dfeovrd(iffcq03aptoverwren),
.ch3_dmonitorclk(iffcq03dmonclk),
.ch3_dmonitorout(iffcq03dmonout),
.ch3_gtrxreset(iffcq03gtrxreset),
.ch3_gttxreset(iffcq03gttxreset),
.ch3_pcsrsvdin(iffcq03pcsrsvdin),
.ch3_phystatus(iffcq03phystatus),
.ch3_rxchbondi(iffcq03rxchbondi),
.ch3_rxchbondo(iffcq03rxchbondo),
.ch3_rxprbserr(iffcq03rxprbserr),
.ch3_rxprbssel(iffcq03rxprbssel),
.ch3_rxqpisenn(iffcq03rxqpisenn),
.ch3_rxqpisenp(iffcq03rxqpisenp),
.ch3_txcominit(iffcq03txcominit),
.ch3_txcomwake(iffcq03txcomwake),
.ch3_txdccdone(iffcq03txdccdone),
.ch3_txdiffctrl(iffcq03txdrvamp),
.ch3_txinhibit(iffcq03txinhibit),
.ch3_txpisopd(iffcq03txserpwrdn),
.ch3_txprbssel(iffcq03txprbssel),
.ch3_txqpisenn(iffcq03txqpisenn),
.ch3_txqpisenp(iffcq03txqpisenp),
.ch3_clkrsvd0(iffcq03ckpinrsrvd0),
.ch3_clkrsvd1(iffcq03ckpinrsrvd1),
.ch3_pinrsvdas(iffcq03pinrsrvdas),
.ch3_rxcdrovrden(iffcq03cdrovren),
.ch3_rxosintdone(iffcq03cfokdone),
.ch3_txprecursor(iffcq03txemppre),
.ch3_cdrstepdir(iffcq03cdrstepdir),
.ch3_pcsrsvdout(iffcq03pcsrsvdout),
.ch3_refdebugout(iffcq03refclkpma),
.ch3_rxcdrreset(iffcq03cdrphreset),
.ch3_rxcommadet(iffcq03rxcommadet),
.ch3_rxcomsasdet(iffcq03comsasdet),
.ch3_rxelecidle(iffcq03rxelecidle),
.ch3_rxoobreset(iffcq03rxoobreset),
.ch3_rxpolarity(iffcq03rxpolarity),
.ch3_rxsliderdy(iffcq03rxsliderdy),
.ch3_rxslipdone(iffcq03rxslipdone),
.ch3_rxsyncdone(iffcq03rxsyncdone),
.ch3_txelecidle(iffcq03txelecidle),
.ch3_txpolarity(iffcq03txpolarity),
.ch3_txpostcursor(iffcq03txemppos),
.ch3_txsequence(iffcq03txsequence),
.ch3_txsyncdone(iffcq03txsyncdone),
.ch3_cdrbmcdrreq(iffcq03cdrbmcdreq),
.ch3_rxclkcorcnt(iffcq03rxckcorcnt),
.ch3_txmaincursor(iffcq03txempmain),
.ch3_bufgtcemask(iffcq03bufgtcemask),
.ch3_cdrincpctrl(iffcq03cdrincpctrl),
.ch3_rxbufstatus(iffcq03rxbufstatus),
.ch3_rxcdrphdone(iffcq03rxcdrphdone),
.ch3_rxcominitdet(iffcq03cominitdet),
.ch3_rxcomwakedet(iffcq03comwakedet),
.ch3_rxdapireset(iffcq03rxdapireset),
.ch3_rxdatavalid(iffcq03rxdatavalid),
.ch3_rxresetdone(iffcq03rxresetdone),
.ch3_rxresetmode(iffcq03rxresetmode),
.ch3_rxsyncallin(iffcq03rxsyncallin),
.ch3_txbufstatus(iffcq03txbufstatus),
.ch3_txcomfinish(iffcq03txcomfinish),
.ch3_txdapireset(iffcq03txdapireset),
.ch3_txoneszeros(iffcq03txoneszeros),
.ch3_txqpibiasen(iffcq03txqpibiasen),
.ch3_txqpiweakpu(iffcq03txqpiweakpu),
.ch3_txresetdone(iffcq03txresetdone),
.ch3_txresetmode(iffcq03txresetmode),
.ch3_txsyncallin(iffcq03txsyncallin),
.ch3_rxphdlypd(iffcq03rxphasealignpd),
.ch3_txphdlypd(iffcq03txphasealignpd),
.ch3_bufgtrstmask(iffcq03bufgtrstmask),
.ch3_eyescanreset(iffcq03eyescanreset),
.ch3_hsdppcsreset(iffcq03hsdppcsreset),
.ch3_iloresetdone(iffcq03iloresetdone),
.ch3_iloresetmask(iffcq03iloresetmask),
.ch3_rxdebugpcsout(iffcq03rxoutpcsclk),
.ch3_rxeqtraining(iffcq03rxeqtraining),
.ch3_rxphdlyreset(iffcq03rxphdlyreset),
.ch3_rxprbslocked(iffcq03rxprbslocked),
.ch3_rxstartofseq(iffcq03rxstartofseq),
.ch3_txdebugpcsout(iffcq03txoutpcsclk),
.ch3_txphdlyreset(iffcq03txphdlyreset),
.ch3_rxmstreset(iffctrlq0mstrxreset[3]),
.ch3_txmstreset(iffctrlq0msttxreset[3]),
.ch3_dmonfiforeset(iffcq03dmonfiforeset),
.ch3_rx10gstat(iffcq03rxethernetstatout),
.ch3_rxbyterealign(q0_ch3_rxbyterealign),
.ch3_rxchanbondseq(iffcq03rxchanbondseq),
.ch3_rxchanrealign(iffcq03rxchanrealign),
.ch3_rxgearboxslip(iffcq03rxgearboxslip),
.ch3_rxheadervalid(iffcq03rxheadervalid),
.ch3_rxmldchainreq(iffcq03rxmldchainreq),
.ch3_rxtermination(iffcq03rxtermination),
.ch3_txmldchainreq(iffcq03txmldchainreq),
.ch3_txpippmstepsize(iffcq03stepsizeppm),
.ch3_txswingoutlow(iffcq03txswingoutlow),
.ch3_rxphalignerr(iffcq03rxphasealignerr),
.ch3_rxphalignreq(iffcq03rxphasealignreq),
.ch3_txphalignerr(iffcq03txphasealignerr),
.ch3_txphalignreq(iffcq03txphasealignreq),
.ch3_txphdlytstclk(iffcq03tcoclkfsmfrout),
.ch3_dmonitoroutclk(q0_ch3_dmonitoroutclk),
.ch3_eyescantrigger(iffcq03eyescantrigger),
.ch3_resetexception(iffcq03resetexception),
.ch3_rxchanisaligned(iffcq03rxchisaligned),
.ch3_rxdlyalignerr(iffcq03rxdelayalignerr),
.ch3_rxdlyalignreq(iffcq03rxdelayalignreq),
.ch3_rxmldchaindone(iffcq03rxmldchaindone),
.ch3_rxpcsresetmask(iffcq03rxpcsresetmask),
.ch3_rxpmaresetdone(iffcq03rxpmaresetdone),
.ch3_rxpmaresetmask(iffcq03rxpmaresetmask),
.ch3_rxprbscntreset(iffcq03rxprbscntreset),
.ch3_rxprogdivreset(iffcq03rxprogdivreset),
.ch3_txdetectrx(iffcq03txdetectrxloopback),
.ch3_txdlyalignerr(iffcq03txdelayalignerr),
.ch3_txdlyalignreq(iffcq03txdelayalignreq),
.ch3_txmldchaindone(iffcq03txmldchaindone),
.ch3_txpcsresetmask(iffcq03txpcsresetmask),
.ch3_txpicodereset(iffcq03txtxpicodereset),
.ch3_txpmaresetdone(iffcq03txpmaresetdone),
.ch3_txpmaresetmask(iffcq03txpmaresetmask),
.ch3_txprbsforceerr(iffcq03txprbsforceerr),
.ch3_txprogdivreset(iffcq03txprogdivreset),
.ch3_txswingouthigh(iffcq03txswingouthigh),
.ch3_rxphaligndone(iffcq03rxphasealigndone),
.ch3_txphaligndone(iffcq03txphasealigndone),
.ch3_rxbyteisaligned(iffcq03rxbyteisaligned),
.ch3_rxdapicodereset(iffcq03rxdapicodereset),
.ch3_rxdapiresetdone(iffcq03rxdapiresetdone),
.ch3_rxdapiresetmask(iffcq03rxdapiresetmask),
.ch3_rxfinealigndone(iffcq03rxfinealigndone),
.ch3_rxphshift180(iffcq03rxphaseshift180req),
.ch3_txdapicodereset(iffcq03txdapicodereset),
.ch3_txdapiresetdone(iffcq03txdapiresetdone),
.ch3_txdapiresetmask(iffcq03txdapiresetmask),
.ch3_txphalignoutrsvd(iffcq03txchicooutrsvd),
.ch3_txphshift180(iffcq03txphaseshift180req),
.ch3_txpicodeovrden(iffcq03txtxpicodeovrden),
.ch3_rxphsetinitreq(iffcq03rxphasesetinitreq),
.ch3_txphsetinitreq(iffcq03txphasesetinitreq),
.ch3_eyescandataerror(iffcq03eyescandataerror),
.ch3_rxdapicodeovrden(iffcq03rxdapicodeovrden),
.ch3_rxmlfinealignreq(iffcq03rxmlfinealignreq),
.ch3_txdapicodeovrden(iffcq03txdapicodeovrden),
.ch3_rxmstresetdone(iffctrlq0mstrxresetdone[3]),
.ch3_rxphsetinitdone(iffcq03rxphasesetinitdone),
.ch3_txmstresetdone(iffctrlq0msttxresetdone[3]),
.ch3_txphsetinitdone(iffcq03txphasesetinitdone),
.ch3_rxdlyalignprog(iffcq03rxdelayalignprogress),
.ch3_rxphalignresetmask(iffcq03rxchicoresetmask),
.ch3_txdlyalignprog(iffcq03txdelayalignprogress),
.ch3_txpausedelayalign(iffcq03txpausedelayalign),
.ch3_txphalignresetmask(iffcq03txchicoresetmask),
.ch3_xpipe5_pipeline_en(iffcq03xpipe5pipelineen),
.ch3_phyesmadaptsave(iffcq03phyesmadaptationsave),
.ch3_rxphshift180done(iffcq03rxphaseshift180done),
.ch3_tx10gstat(iffcq03txethernetstattxlocalfault),
.ch3_txphshift180done(iffcq03txphaseshift180done),
.ch3_rxprogdivresetdone(iffcq03rxprogdivresetdone),
.ch3_rxsimplexphystatus(iffcq03rxsimplexphystatus),
.ch3_txprogdivresetdone(iffcq03txprogdivresetdone),
.ch3_txsimplexphystatus(iffcq03txsimplexphystatus),
.ch3_rxphdlyresetdone(iffcq03rxphasedelayresetdone),
.ch3_txphdlyresetdone(iffcq03txphasedelayresetdone),

.ctrlrsvdin(iffctrlq0gtrsvdin),
.ctrlrsvdout(iffctrlq0gtrsvdout),
.coestatusdebug(iffctrlq0coeregrst),
.correcterr(iffctrlq0correctableerr),

.debugtraceclk(iffctrlq0debugtraceclk),
.debugtracetdata(iffctrlq0debugtracetdata),
.debugtraceready(iffctrlq0debugtracetready),
.debugtracetvalid(iffctrlq0debugtracetvalid),

.gpi(iffctrlq0ubgpi),
.gpo(iffctrlq0ubgpo),
.gtpowergood(iffctrlq0gtpowergood),

.hsclk0_rpllpd(iffhsq00rpllpwrdn),
.hsclk0_lcpllpd(iffhsq00lcpllpwrdn),
.hsclk0_rpllfbdiv(iffhsq00rpllfbdiv),
.hsclk0_rpllreset(iffhsq00rpllreset),
.hsclk0_lcpllfbdiv(iffhsq00lcpllfbdiv),
.hsclk0_lcpllreset(iffhsq00lcpllreset),
.hsclk0_rplllock(iffhsq00rpllfreqlock),
.hsclk0_lcplllock(iffhsq00lcpllfreqlock),
.hsclk0_rpllsdmdata(iffhsq00rpllsdmdata),
.hsclk0_rpllfbclklost(iffhsq00rpllfbloss),
.hsclk0_lcpllsdmdata(iffhsq00lcpllsdmdata),
.hsclk0_rxrecclkout0(iffhsq00rxrecclkout0),
.hsclk0_rxrecclkout1(iffhsq00rxrecclkout1),
.hsclk0_lcpllfbclklost(iffhsq00lcpllfbloss),
.hsclk0_rpllrefclklost(iffhsq00rpllrefloss),
.hsclk0_rpllrefclksel(iffhsq00rpllrefseldyn),
.hsclk0_rpllresetmask(iffhsq00rpllresetmask),
.hsclk0_rpllsdmtoggle(iffhsq00rpllsdmtoggle),
.hsclk0_lcpllrefclklost(iffhsq00lcpllrefloss),
.hsclk0_lcpllrefclksel(iffhsq00lcpllrefseldyn),
.hsclk0_lcpllresetmask(iffhsq00lcpllresetmask),
.hsclk0_lcpllsdmtoggle(iffhsq00lcpllsdmtoggle),
.hsclk0_rpllrefclkmonitor(iffhsq00mgtrpllrefclkfa),
.hsclk0_lcpllrefclkmonitor(iffhsq00mgtlcpllrefclkfa),
.hsclk0_rpllresetbypassmode(iffhsq00rpllresetbypassmode),
.hsclk0_lcpllresetbypassmode(iffhsq00lcpllresetbypassmode),

.hsclk1_rpllpd(iffhsq01rpllpwrdn),
.hsclk1_lcpllpd(iffhsq01lcpllpwrdn),
.hsclk1_rpllfbdiv(iffhsq01rpllfbdiv),
.hsclk1_rpllreset(iffhsq01rpllreset),
.hsclk1_lcpllfbdiv(iffhsq01lcpllfbdiv),
.hsclk1_lcpllreset(iffhsq01lcpllreset),
.hsclk1_rplllock(iffhsq01rpllfreqlock),
.hsclk1_lcplllock(iffhsq01lcpllfreqlock),
.hsclk1_rpllsdmdata(iffhsq01rpllsdmdata),
.hsclk1_rpllfbclklost(iffhsq01rpllfbloss),
.hsclk1_lcpllsdmdata(iffhsq01lcpllsdmdata),
.hsclk1_rxrecclkout0(iffhsq01rxrecclkout0),
.hsclk1_rxrecclkout1(iffhsq01rxrecclkout1),
.hsclk1_lcpllfbclklost(iffhsq01lcpllfbloss),
.hsclk1_rpllrefclklost(iffhsq01rpllrefloss),
.hsclk1_rpllrefclksel(iffhsq01rpllrefseldyn),
.hsclk1_rpllresetmask(iffhsq01rpllresetmask),
.hsclk1_rpllsdmtoggle(iffhsq01rpllsdmtoggle),
.hsclk1_lcpllrefclklost(iffhsq01lcpllrefloss),
.hsclk1_lcpllrefclksel(iffhsq01lcpllrefseldyn),
.hsclk1_lcpllresetmask(iffhsq01lcpllresetmask),
.hsclk1_lcpllsdmtoggle(iffhsq01lcpllsdmtoggle),
.hsclk1_rpllrefclkmonitor(iffhsq01mgtrpllrefclkfa),
.hsclk1_lcpllrefclkmonitor(iffhsq01mgtlcpllrefclkfa),
.hsclk1_rpllresetbypassmode(iffhsq01rpllresetbypassmode),
.hsclk1_lcpllresetbypassmode(iffhsq01lcpllresetbypassmode),

.m0_axis_tdata(iffctrlq0m0axistdata),
.m0_axis_tlast(iffctrlq0m0axistlast),
.m1_axis_tdata(iffctrlq0m1axistdata),
.m1_axis_tlast(iffctrlq0m1axistlast),
.m2_axis_tdata(iffctrlq0m2axistdata),
.m2_axis_tlast(iffctrlq0m2axistlast),
.s0_axis_tdata(iffctrlq0s0axistdata),
.s0_axis_tlast(iffctrlq0s0axistlast),
.s1_axis_tdata(iffctrlq0s1axistdata),
.s1_axis_tlast(iffctrlq0s1axistlast),
.s2_axis_tdata(iffctrlq0s2axistdata),
.s2_axis_tlast(iffctrlq0s2axistlast),
.m0_axis_tready(iffctrlq0m0axistready),
.m0_axis_tvalid(iffctrlq0m0axistvalid),
.m1_axis_tready(iffctrlq0m1axistready),
.m1_axis_tvalid(iffctrlq0m1axistvalid),
.m2_axis_tready(iffctrlq0m2axistready),
.m2_axis_tvalid(iffctrlq0m2axistvalid),
.s0_axis_tready(iffctrlq0s0axistready),
.s0_axis_tvalid(iffctrlq0s0axistvalid),
.s1_axis_tready(iffctrlq0s1axistready),
.s1_axis_tvalid(iffctrlq0s1axistvalid),
.s2_axis_tready(iffctrlq0s2axistready),
.s2_axis_tvalid(iffctrlq0s2axistvalid),

.rcalenb(iffctrlq0rcalenb),
.pcieltssm(iffctrlq0pcieltssmstate),
.uncorrecterr(iffctrlq0uncorrectableerr),
.pcielinkreachtarget(iffctrlq0pcielinkreachtarget),

.refclk0_clktestsigint(),
.refclk1_clktestsigint(),
.refclk0_gtrefclkpd(iffrckq00refclkpd),
.refclk1_gtrefclkpd(iffrckq01refclkpd),
.refclk0_clktestsig(iffrckq00hrowtestck),
.refclk1_clktestsig(iffrckq01hrowtestck),
.refclk0_gtrefclkpdint(gt0_refclk0_pdint),
.refclk1_gtrefclkpdint(gt0_refclk1_pdint),

.rxmarginclk(iffctrlq0rxmarginclk),
.rxmarginreqack(iffctrlq0rxmarginreqack),
.rxmarginreqcmd(iffctrlq0rxmarginreqcmd),
.rxmarginreqreq(iffctrlq0rxmarginreqreq),
.rxmarginresack(iffctrlq0rxmarginresack),
.rxmarginrescmd(iffctrlq0rxmarginrescmd),
.rxmarginresreq(iffctrlq0rxmarginresreq),
.rxmarginrespayld(iffctrlq0rxmarginrespayld),
.rxmarginreqpayld(iffctrlq0rxmarginreqpayload),
.rxmarginreqlanenum(iffctrlq0rxmarginreqlanenum),
.rxmarginreslanenum(iffctrlq0rxmarginreslanenum),

.trigin0(iffctrlq0trigin0),
.trigout0(iffctrlq0trigout0),
.trigackin0(iffctrlq0trigackin0),
.trigackout0(iffctrlq0trigackout0),

.ubintr(iffctrlq0ubintr),
.ubmbrst(iffctrlq0ubmbrst),
.ubenable(iffctrlq0ubenable),
.ubrxuart(iffctrlq0ubrxuart),
.ubtxuart(iffctrlq0ubtxuart),
.ubiolmbrst(iffctrlq0ubiolmbrst),
.ubinterrupt(iffctrlq0ubinterrupt),

.pipesouthout(),
.rxpisouthout(),
.txpisouthout(),
.pipenorthin('d0),
.rxpinorthin('d0),
.txpinorthin('d0),
.resetdone_southout(),
.resetdone_northin('d0),
.rxpisouthin(rxpisouthin_to_rxpsouthout_q1),
.txpisouthin(txpisouthin_to_txpsouthout_q1),
.pipenorthout(pipenorthoutq0_to_pipenorthinq1),
.pipesouthin(pipesouthin_q0_to_pipesouthout_q1),
.rxpinorthout(rxpinorthout_q0_to_rxpinorthin_q1),
.txpinorthout(txpinorthout_q0_to_txpinorthin_q1),
.resetdone_southin(resetdone_southin_q0_to_resetdone_southout_q1),
.resetdone_northout(resetdone_northout_q0_to_resetdone_northin_q1),

.rxn(gt0_serial_rxn),
.rxp(gt0_serial_rxp),
.txn(gt0_serial_txn),
.txp(gt0_serial_txp)
